magic
tech sky130A
magscale 1 2
timestamp 1740018547
<< viali >>
rect 8033 18921 8067 18955
rect 8677 18921 8711 18955
rect 9965 18921 9999 18955
rect 10609 18921 10643 18955
rect 11253 18921 11287 18955
rect 13829 18921 13863 18955
rect 7849 18717 7883 18751
rect 8493 18717 8527 18751
rect 9781 18717 9815 18751
rect 10425 18717 10459 18751
rect 11069 18717 11103 18751
rect 13645 18717 13679 18751
rect 14473 18717 14507 18751
rect 13461 18649 13495 18683
rect 14749 18649 14783 18683
rect 13369 18581 13403 18615
rect 16221 18581 16255 18615
rect 7573 18377 7607 18411
rect 10057 18377 10091 18411
rect 11253 18377 11287 18411
rect 12357 18377 12391 18411
rect 13369 18377 13403 18411
rect 10793 18309 10827 18343
rect 14289 18309 14323 18343
rect 7941 18241 7975 18275
rect 8033 18241 8067 18275
rect 8401 18241 8435 18275
rect 8585 18241 8619 18275
rect 8861 18241 8895 18275
rect 8953 18241 8987 18275
rect 9137 18241 9171 18275
rect 9229 18241 9263 18275
rect 9413 18241 9447 18275
rect 9505 18241 9539 18275
rect 9873 18241 9907 18275
rect 10885 18241 10919 18275
rect 11529 18241 11563 18275
rect 11713 18241 11747 18275
rect 12081 18241 12115 18275
rect 13001 18241 13035 18275
rect 13553 18241 13587 18275
rect 13645 18241 13679 18275
rect 16037 18241 16071 18275
rect 8125 18173 8159 18207
rect 8769 18173 8803 18207
rect 9689 18173 9723 18207
rect 10701 18173 10735 18207
rect 11989 18173 12023 18207
rect 12357 18173 12391 18207
rect 13093 18173 13127 18207
rect 14013 18173 14047 18207
rect 9137 18105 9171 18139
rect 9229 18105 9263 18139
rect 15761 18105 15795 18139
rect 11897 18037 11931 18071
rect 12173 18037 12207 18071
rect 13829 18037 13863 18071
rect 15945 18037 15979 18071
rect 9689 17833 9723 17867
rect 10057 17833 10091 17867
rect 10701 17833 10735 17867
rect 11989 17833 12023 17867
rect 12357 17833 12391 17867
rect 13461 17833 13495 17867
rect 16681 17833 16715 17867
rect 11805 17765 11839 17799
rect 9965 17697 9999 17731
rect 12081 17697 12115 17731
rect 13277 17697 13311 17731
rect 14749 17697 14783 17731
rect 2605 17629 2639 17663
rect 10057 17629 10091 17663
rect 11529 17629 11563 17663
rect 11805 17629 11839 17663
rect 11989 17629 12023 17663
rect 13185 17629 13219 17663
rect 14473 17629 14507 17663
rect 16773 17629 16807 17663
rect 10333 17561 10367 17595
rect 10517 17561 10551 17595
rect 16497 17561 16531 17595
rect 2697 17493 2731 17527
rect 11621 17493 11655 17527
rect 5733 17289 5767 17323
rect 7021 17289 7055 17323
rect 10425 17289 10459 17323
rect 10885 17289 10919 17323
rect 13737 17289 13771 17323
rect 14197 17289 14231 17323
rect 9045 17221 9079 17255
rect 10057 17221 10091 17255
rect 11069 17221 11103 17255
rect 16773 17221 16807 17255
rect 3893 17153 3927 17187
rect 3985 17153 4019 17187
rect 5365 17153 5399 17187
rect 5825 17153 5859 17187
rect 5917 17153 5951 17187
rect 6561 17153 6595 17187
rect 6837 17153 6871 17187
rect 7297 17153 7331 17187
rect 8033 17153 8067 17187
rect 8585 17153 8619 17187
rect 8677 17153 8711 17187
rect 8953 17153 8987 17187
rect 9505 17153 9539 17187
rect 9873 17153 9907 17187
rect 10149 17153 10183 17187
rect 10241 17153 10275 17187
rect 10609 17153 10643 17187
rect 11253 17153 11287 17187
rect 11805 17153 11839 17187
rect 12265 17153 12299 17187
rect 13369 17153 13403 17187
rect 13829 17153 13863 17187
rect 14013 17153 14047 17187
rect 16497 17153 16531 17187
rect 4169 17085 4203 17119
rect 7665 17085 7699 17119
rect 9229 17085 9263 17119
rect 9781 17085 9815 17119
rect 11529 17085 11563 17119
rect 13277 17085 13311 17119
rect 13461 17085 13495 17119
rect 13553 17085 13587 17119
rect 14749 17085 14783 17119
rect 6009 17017 6043 17051
rect 8401 16949 8435 16983
rect 10701 16949 10735 16983
rect 16865 16949 16899 16983
rect 7665 16745 7699 16779
rect 10333 16745 10367 16779
rect 13737 16745 13771 16779
rect 15117 16745 15151 16779
rect 5181 16677 5215 16711
rect 13093 16677 13127 16711
rect 3617 16609 3651 16643
rect 3985 16609 4019 16643
rect 4077 16609 4111 16643
rect 4169 16609 4203 16643
rect 4537 16609 4571 16643
rect 5365 16609 5399 16643
rect 5549 16609 5583 16643
rect 7205 16609 7239 16643
rect 7757 16609 7791 16643
rect 7941 16609 7975 16643
rect 8033 16609 8067 16643
rect 8217 16609 8251 16643
rect 10149 16609 10183 16643
rect 14933 16609 14967 16643
rect 3249 16541 3283 16575
rect 3433 16541 3467 16575
rect 4261 16541 4295 16575
rect 4721 16541 4755 16575
rect 4813 16541 4847 16575
rect 4997 16541 5031 16575
rect 5089 16541 5123 16575
rect 5457 16541 5491 16575
rect 5641 16541 5675 16575
rect 6101 16541 6135 16575
rect 6929 16541 6963 16575
rect 7113 16541 7147 16575
rect 7297 16541 7331 16575
rect 7481 16541 7515 16575
rect 8125 16541 8159 16575
rect 8769 16541 8803 16575
rect 8953 16541 8987 16575
rect 9873 16541 9907 16575
rect 10241 16541 10275 16575
rect 10425 16541 10459 16575
rect 10793 16541 10827 16575
rect 11069 16541 11103 16575
rect 12909 16541 12943 16575
rect 13093 16541 13127 16575
rect 13277 16541 13311 16575
rect 13645 16541 13679 16575
rect 13829 16541 13863 16575
rect 15025 16541 15059 16575
rect 15761 16541 15795 16575
rect 16221 16541 16255 16575
rect 16497 16541 16531 16575
rect 16589 16541 16623 16575
rect 6469 16473 6503 16507
rect 6653 16473 6687 16507
rect 15853 16473 15887 16507
rect 4445 16405 4479 16439
rect 5917 16405 5951 16439
rect 6837 16405 6871 16439
rect 8585 16405 8619 16439
rect 9137 16405 9171 16439
rect 10609 16405 10643 16439
rect 13461 16405 13495 16439
rect 14703 16405 14737 16439
rect 5641 16201 5675 16235
rect 6929 16201 6963 16235
rect 7665 16201 7699 16235
rect 8309 16201 8343 16235
rect 8677 16201 8711 16235
rect 11161 16201 11195 16235
rect 15853 16201 15887 16235
rect 6529 16133 6563 16167
rect 6745 16133 6779 16167
rect 8125 16133 8159 16167
rect 9873 16133 9907 16167
rect 11897 16133 11931 16167
rect 12081 16133 12115 16167
rect 12265 16133 12299 16167
rect 12449 16133 12483 16167
rect 12909 16133 12943 16167
rect 13093 16133 13127 16167
rect 13553 16133 13587 16167
rect 16037 16133 16071 16167
rect 17141 16133 17175 16167
rect 2789 16065 2823 16099
rect 3157 16065 3191 16099
rect 5641 16065 5675 16099
rect 6101 16065 6135 16099
rect 6837 16065 6871 16099
rect 7113 16065 7147 16099
rect 7205 16065 7239 16099
rect 7389 16065 7423 16099
rect 7481 16065 7515 16099
rect 7941 16065 7975 16099
rect 8585 16065 8619 16099
rect 8861 16065 8895 16099
rect 9321 16065 9355 16099
rect 10057 16065 10091 16099
rect 10701 16065 10735 16099
rect 11069 16065 11103 16099
rect 11253 16065 11287 16099
rect 11529 16065 11563 16099
rect 11713 16065 11747 16099
rect 11805 16065 11839 16099
rect 11989 16065 12023 16099
rect 12725 16065 12759 16099
rect 12817 16065 12851 16099
rect 13369 16065 13403 16099
rect 13829 16065 13863 16099
rect 14105 16065 14139 16099
rect 16129 16065 16163 16099
rect 16865 16065 16899 16099
rect 5089 15997 5123 16031
rect 5181 15997 5215 16031
rect 5273 15997 5307 16031
rect 5365 15997 5399 16031
rect 5549 15997 5583 16031
rect 5825 15997 5859 16031
rect 7297 15997 7331 16031
rect 9597 15997 9631 16031
rect 10241 15997 10275 16031
rect 10977 15997 11011 16031
rect 13185 15997 13219 16031
rect 13645 15997 13679 16031
rect 14013 15997 14047 16031
rect 14381 15997 14415 16031
rect 5963 15929 5997 15963
rect 7113 15929 7147 15963
rect 10793 15929 10827 15963
rect 12541 15929 12575 15963
rect 4445 15861 4479 15895
rect 6377 15861 6411 15895
rect 6561 15861 6595 15895
rect 9045 15861 9079 15895
rect 10885 15861 10919 15895
rect 11621 15861 11655 15895
rect 16773 15861 16807 15895
rect 17233 15861 17267 15895
rect 2697 15657 2731 15691
rect 3249 15657 3283 15691
rect 4537 15657 4571 15691
rect 9965 15657 9999 15691
rect 15117 15657 15151 15691
rect 2881 15589 2915 15623
rect 9137 15589 9171 15623
rect 4445 15521 4479 15555
rect 4997 15521 5031 15555
rect 8585 15521 8619 15555
rect 9045 15521 9079 15555
rect 15301 15521 15335 15555
rect 17233 15521 17267 15555
rect 2513 15453 2547 15487
rect 2697 15453 2731 15487
rect 4261 15453 4295 15487
rect 4905 15453 4939 15487
rect 5181 15453 5215 15487
rect 5273 15453 5307 15487
rect 5549 15453 5583 15487
rect 5917 15453 5951 15487
rect 6469 15453 6503 15487
rect 7757 15453 7791 15487
rect 7905 15453 7939 15487
rect 8125 15453 8159 15487
rect 8222 15453 8256 15487
rect 8677 15453 8711 15487
rect 9413 15453 9447 15487
rect 9505 15453 9539 15487
rect 9873 15453 9907 15487
rect 9965 15453 9999 15487
rect 12725 15453 12759 15487
rect 14933 15453 14967 15487
rect 17141 15453 17175 15487
rect 17543 15453 17577 15487
rect 3249 15385 3283 15419
rect 4537 15385 4571 15419
rect 5457 15385 5491 15419
rect 6653 15385 6687 15419
rect 8033 15385 8067 15419
rect 9321 15385 9355 15419
rect 15577 15385 15611 15419
rect 3433 15317 3467 15351
rect 4077 15317 4111 15351
rect 8401 15317 8435 15351
rect 9781 15317 9815 15351
rect 10241 15317 10275 15351
rect 12909 15317 12943 15351
rect 17049 15317 17083 15351
rect 17693 15317 17727 15351
rect 7757 15113 7791 15147
rect 8861 15113 8895 15147
rect 11529 15113 11563 15147
rect 12357 15113 12391 15147
rect 15209 15113 15243 15147
rect 16865 15113 16899 15147
rect 17693 15113 17727 15147
rect 3801 15045 3835 15079
rect 7297 15045 7331 15079
rect 9397 15045 9431 15079
rect 9597 15045 9631 15079
rect 10701 15045 10735 15079
rect 10793 15045 10827 15079
rect 12725 15045 12759 15079
rect 12843 15045 12877 15079
rect 16497 15045 16531 15079
rect 2053 14977 2087 15011
rect 2329 14977 2363 15011
rect 2421 14977 2455 15011
rect 2605 14977 2639 15011
rect 2697 14977 2731 15011
rect 3065 14977 3099 15011
rect 3985 14977 4019 15011
rect 4169 14977 4203 15011
rect 4261 14977 4295 15011
rect 5549 14977 5583 15011
rect 5733 14977 5767 15011
rect 7205 14977 7239 15011
rect 7389 14977 7423 15011
rect 7573 14977 7607 15011
rect 7665 14977 7699 15011
rect 7941 14977 7975 15011
rect 9045 14977 9079 15011
rect 9965 14977 9999 15011
rect 10425 14977 10459 15011
rect 10517 14977 10551 15011
rect 10885 14977 10919 15011
rect 12081 14977 12115 15011
rect 12541 14977 12575 15011
rect 12633 14977 12667 15011
rect 13369 14977 13403 15011
rect 13461 14977 13495 15011
rect 16681 14977 16715 15011
rect 16957 14977 16991 15011
rect 17049 14977 17083 15011
rect 17969 14977 18003 15011
rect 1777 14909 1811 14943
rect 2145 14909 2179 14943
rect 2789 14909 2823 14943
rect 2973 14909 3007 14943
rect 3157 14909 3191 14943
rect 3249 14909 3283 14943
rect 8125 14909 8159 14943
rect 11805 14909 11839 14943
rect 13001 14909 13035 14943
rect 13277 14909 13311 14943
rect 13553 14909 13587 14943
rect 9781 14841 9815 14875
rect 11069 14841 11103 14875
rect 17233 14841 17267 14875
rect 1869 14773 1903 14807
rect 1961 14773 1995 14807
rect 5917 14773 5951 14807
rect 7021 14773 7055 14807
rect 9229 14773 9263 14807
rect 9413 14773 9447 14807
rect 11713 14773 11747 14807
rect 13093 14773 13127 14807
rect 16681 14773 16715 14807
rect 2329 14569 2363 14603
rect 6377 14569 6411 14603
rect 6469 14569 6503 14603
rect 7205 14569 7239 14603
rect 9321 14569 9355 14603
rect 10241 14569 10275 14603
rect 11805 14569 11839 14603
rect 12817 14569 12851 14603
rect 1501 14501 1535 14535
rect 7297 14501 7331 14535
rect 10885 14501 10919 14535
rect 14105 14501 14139 14535
rect 16313 14501 16347 14535
rect 6285 14433 6319 14467
rect 7573 14433 7607 14467
rect 7757 14433 7791 14467
rect 8677 14433 8711 14467
rect 9229 14433 9263 14467
rect 12725 14433 12759 14467
rect 15669 14433 15703 14467
rect 15761 14433 15795 14467
rect 16129 14433 16163 14467
rect 18061 14433 18095 14467
rect 1685 14365 1719 14399
rect 2329 14365 2363 14399
rect 2513 14365 2547 14399
rect 2605 14365 2639 14399
rect 4169 14365 4203 14399
rect 4353 14365 4387 14399
rect 4445 14365 4479 14399
rect 4721 14365 4755 14399
rect 4905 14365 4939 14399
rect 4997 14365 5031 14399
rect 6193 14365 6227 14399
rect 6561 14365 6595 14399
rect 6653 14365 6687 14399
rect 7021 14365 7055 14399
rect 7481 14365 7515 14399
rect 7665 14365 7699 14399
rect 8585 14365 8619 14399
rect 8769 14365 8803 14399
rect 8953 14365 8987 14399
rect 9597 14365 9631 14399
rect 9781 14365 9815 14399
rect 9873 14365 9907 14399
rect 9965 14365 9999 14399
rect 10793 14365 10827 14399
rect 10977 14365 11011 14399
rect 11161 14365 11195 14399
rect 11309 14365 11343 14399
rect 11645 14365 11679 14399
rect 12357 14365 12391 14399
rect 12541 14365 12575 14399
rect 12633 14365 12667 14399
rect 14289 14365 14323 14399
rect 14657 14365 14691 14399
rect 14749 14365 14783 14399
rect 14841 14365 14875 14399
rect 14933 14365 14967 14399
rect 15301 14365 15335 14399
rect 15853 14365 15887 14399
rect 15945 14365 15979 14399
rect 5917 14297 5951 14331
rect 6837 14297 6871 14331
rect 6929 14297 6963 14331
rect 11437 14297 11471 14331
rect 11529 14297 11563 14331
rect 12909 14297 12943 14331
rect 14381 14297 14415 14331
rect 14473 14297 14507 14331
rect 15117 14297 15151 14331
rect 15209 14297 15243 14331
rect 17785 14297 17819 14331
rect 3985 14229 4019 14263
rect 4537 14229 4571 14263
rect 5181 14229 5215 14263
rect 9505 14229 9539 14263
rect 15485 14229 15519 14263
rect 2697 14025 2731 14059
rect 4169 14025 4203 14059
rect 6009 14025 6043 14059
rect 9505 14025 9539 14059
rect 11529 14025 11563 14059
rect 14749 14025 14783 14059
rect 16957 14025 16991 14059
rect 17049 14025 17083 14059
rect 17509 14025 17543 14059
rect 17969 14025 18003 14059
rect 3249 13957 3283 13991
rect 5549 13957 5583 13991
rect 5749 13957 5783 13991
rect 1685 13889 1719 13923
rect 2513 13889 2547 13923
rect 2789 13889 2823 13923
rect 3065 13889 3099 13923
rect 3893 13889 3927 13923
rect 5181 13889 5215 13923
rect 5273 13889 5307 13923
rect 5365 13889 5399 13923
rect 6009 13889 6043 13923
rect 6193 13889 6227 13923
rect 6929 13889 6963 13923
rect 7113 13889 7147 13923
rect 7389 13889 7423 13923
rect 7573 13889 7607 13923
rect 7941 13889 7975 13923
rect 8033 13889 8067 13923
rect 8217 13889 8251 13923
rect 8309 13889 8343 13923
rect 8585 13889 8619 13923
rect 8861 13889 8895 13923
rect 8953 13889 8987 13923
rect 9413 13889 9447 13923
rect 9597 13889 9631 13923
rect 10057 13889 10091 13923
rect 11069 13889 11103 13923
rect 11253 13889 11287 13923
rect 11345 13911 11379 13945
rect 11713 13889 11747 13923
rect 11805 13889 11839 13923
rect 14289 13889 14323 13923
rect 14381 13889 14415 13923
rect 14657 13889 14691 13923
rect 14933 13889 14967 13923
rect 15025 13889 15059 13923
rect 16221 13889 16255 13923
rect 16681 13889 16715 13923
rect 17049 13889 17083 13923
rect 17233 13889 17267 13923
rect 17325 13889 17359 13923
rect 17509 13889 17543 13923
rect 17785 13889 17819 13923
rect 4169 13821 4203 13855
rect 7205 13821 7239 13855
rect 7297 13821 7331 13855
rect 12173 13821 12207 13855
rect 14105 13821 14139 13855
rect 14197 13821 14231 13855
rect 14565 13821 14599 13855
rect 14841 13821 14875 13855
rect 15669 13821 15703 13855
rect 15945 13821 15979 13855
rect 16037 13821 16071 13855
rect 16957 13821 16991 13855
rect 5917 13753 5951 13787
rect 8493 13753 8527 13787
rect 1501 13685 1535 13719
rect 2329 13685 2363 13719
rect 2881 13685 2915 13719
rect 3985 13685 4019 13719
rect 5724 13685 5758 13719
rect 8677 13685 8711 13719
rect 9137 13685 9171 13719
rect 9781 13685 9815 13719
rect 10885 13685 10919 13719
rect 16773 13685 16807 13719
rect 3341 13481 3375 13515
rect 4169 13481 4203 13515
rect 7113 13481 7147 13515
rect 7297 13481 7331 13515
rect 8953 13481 8987 13515
rect 10793 13481 10827 13515
rect 13185 13481 13219 13515
rect 15393 13481 15427 13515
rect 16037 13481 16071 13515
rect 17785 13481 17819 13515
rect 1777 13413 1811 13447
rect 2605 13413 2639 13447
rect 8677 13413 8711 13447
rect 12817 13413 12851 13447
rect 2053 13345 2087 13379
rect 9137 13345 9171 13379
rect 9597 13345 9631 13379
rect 9689 13345 9723 13379
rect 9873 13345 9907 13379
rect 10517 13345 10551 13379
rect 11161 13345 11195 13379
rect 11253 13345 11287 13379
rect 1501 13277 1535 13311
rect 1593 13277 1627 13311
rect 1777 13277 1811 13311
rect 2976 13277 3010 13311
rect 3157 13277 3191 13311
rect 3801 13277 3835 13311
rect 3985 13277 4019 13311
rect 5273 13277 5307 13311
rect 5457 13277 5491 13311
rect 7389 13277 7423 13311
rect 7665 13277 7699 13311
rect 8585 13277 8619 13311
rect 8769 13277 8803 13311
rect 9229 13277 9263 13311
rect 9965 13277 9999 13311
rect 10057 13277 10091 13311
rect 10149 13277 10183 13311
rect 10425 13277 10459 13311
rect 10609 13277 10643 13311
rect 10977 13277 11011 13311
rect 11069 13277 11103 13311
rect 13001 13277 13035 13311
rect 13277 13277 13311 13311
rect 13369 13277 13403 13311
rect 13553 13277 13587 13311
rect 14933 13277 14967 13311
rect 15209 13277 15243 13311
rect 15853 13277 15887 13311
rect 2605 13209 2639 13243
rect 3433 13209 3467 13243
rect 5365 13209 5399 13243
rect 9505 13209 9539 13243
rect 16313 13209 16347 13243
rect 1869 13141 1903 13175
rect 2145 13141 2179 13175
rect 2789 13141 2823 13175
rect 13553 13141 13587 13175
rect 15025 13141 15059 13175
rect 1501 12937 1535 12971
rect 1961 12937 1995 12971
rect 2605 12937 2639 12971
rect 3617 12937 3651 12971
rect 6377 12937 6411 12971
rect 15945 12937 15979 12971
rect 17785 12937 17819 12971
rect 1869 12869 1903 12903
rect 2973 12869 3007 12903
rect 5733 12869 5767 12903
rect 6863 12869 6897 12903
rect 9045 12869 9079 12903
rect 11529 12869 11563 12903
rect 14657 12869 14691 12903
rect 14841 12869 14875 12903
rect 2789 12801 2823 12835
rect 3065 12801 3099 12835
rect 3801 12801 3835 12835
rect 3893 12801 3927 12835
rect 4077 12801 4111 12835
rect 4261 12801 4295 12835
rect 4721 12801 4755 12835
rect 4905 12801 4939 12835
rect 5089 12801 5123 12835
rect 5917 12801 5951 12835
rect 6101 12801 6135 12835
rect 6561 12801 6595 12835
rect 6653 12801 6687 12835
rect 6745 12801 6779 12835
rect 7021 12801 7055 12835
rect 8953 12801 8987 12835
rect 9137 12801 9171 12835
rect 9781 12801 9815 12835
rect 9873 12801 9907 12835
rect 10793 12801 10827 12835
rect 11805 12801 11839 12835
rect 11897 12801 11931 12835
rect 11989 12801 12023 12835
rect 13093 12801 13127 12835
rect 13277 12801 13311 12835
rect 13645 12801 13679 12835
rect 13737 12801 13771 12835
rect 14197 12801 14231 12835
rect 14381 12801 14415 12835
rect 14933 12801 14967 12835
rect 15301 12801 15335 12835
rect 15577 12801 15611 12835
rect 15853 12801 15887 12835
rect 16129 12801 16163 12835
rect 16497 12801 16531 12835
rect 16681 12801 16715 12835
rect 17325 12801 17359 12835
rect 17601 12801 17635 12835
rect 17693 12801 17727 12835
rect 2053 12733 2087 12767
rect 3985 12733 4019 12767
rect 4997 12733 5031 12767
rect 6193 12733 6227 12767
rect 9689 12733 9723 12767
rect 9965 12733 9999 12767
rect 10701 12733 10735 12767
rect 11529 12733 11563 12767
rect 12173 12733 12207 12767
rect 13461 12733 13495 12767
rect 13553 12733 13587 12767
rect 15117 12733 15151 12767
rect 10425 12665 10459 12699
rect 11897 12665 11931 12699
rect 14289 12665 14323 12699
rect 15025 12665 15059 12699
rect 17233 12665 17267 12699
rect 4629 12597 4663 12631
rect 9505 12597 9539 12631
rect 10793 12597 10827 12631
rect 11713 12597 11747 12631
rect 13185 12597 13219 12631
rect 13921 12597 13955 12631
rect 14657 12597 14691 12631
rect 16129 12597 16163 12631
rect 16865 12597 16899 12631
rect 17509 12597 17543 12631
rect 2421 12393 2455 12427
rect 3985 12393 4019 12427
rect 4261 12393 4295 12427
rect 6745 12393 6779 12427
rect 7757 12393 7791 12427
rect 8585 12393 8619 12427
rect 9597 12393 9631 12427
rect 11253 12393 11287 12427
rect 11345 12393 11379 12427
rect 11805 12393 11839 12427
rect 12909 12393 12943 12427
rect 15577 12393 15611 12427
rect 15945 12393 15979 12427
rect 5733 12325 5767 12359
rect 6929 12325 6963 12359
rect 5825 12257 5859 12291
rect 6653 12257 6687 12291
rect 11437 12257 11471 12291
rect 13461 12257 13495 12291
rect 2605 12189 2639 12223
rect 2973 12189 3007 12223
rect 3065 12189 3099 12223
rect 4445 12189 4479 12223
rect 4813 12189 4847 12223
rect 4905 12189 4939 12223
rect 5273 12189 5307 12223
rect 5457 12189 5491 12223
rect 6561 12189 6595 12223
rect 7205 12189 7239 12223
rect 7297 12189 7331 12223
rect 7389 12189 7423 12223
rect 7481 12189 7515 12223
rect 7665 12189 7699 12223
rect 7941 12189 7975 12223
rect 8309 12189 8343 12223
rect 9137 12189 9171 12223
rect 9321 12189 9355 12223
rect 11069 12189 11103 12223
rect 11253 12189 11287 12223
rect 11621 12189 11655 12223
rect 11897 12189 11931 12223
rect 12081 12189 12115 12223
rect 12633 12189 12667 12223
rect 12725 12189 12759 12223
rect 12909 12189 12943 12223
rect 13185 12189 13219 12223
rect 13369 12189 13403 12223
rect 13553 12189 13587 12223
rect 13737 12189 13771 12223
rect 14381 12189 14415 12223
rect 14473 12189 14507 12223
rect 14657 12189 14691 12223
rect 14749 12189 14783 12223
rect 15117 12189 15151 12223
rect 15485 12189 15519 12223
rect 15669 12189 15703 12223
rect 17693 12189 17727 12223
rect 2697 12121 2731 12155
rect 2789 12121 2823 12155
rect 3801 12121 3835 12155
rect 4537 12121 4571 12155
rect 4629 12121 4663 12155
rect 8585 12121 8619 12155
rect 9689 12121 9723 12155
rect 11345 12121 11379 12155
rect 17417 12121 17451 12155
rect 4001 12053 4035 12087
rect 4169 12053 4203 12087
rect 7021 12053 7055 12087
rect 8217 12053 8251 12087
rect 8401 12053 8435 12087
rect 9137 12053 9171 12087
rect 12081 12053 12115 12087
rect 13001 12053 13035 12087
rect 14933 12053 14967 12087
rect 15301 12053 15335 12087
rect 3065 11849 3099 11883
rect 4353 11849 4387 11883
rect 7205 11849 7239 11883
rect 7849 11849 7883 11883
rect 13001 11849 13035 11883
rect 3985 11781 4019 11815
rect 7665 11781 7699 11815
rect 9597 11781 9631 11815
rect 9689 11781 9723 11815
rect 2421 11713 2455 11747
rect 2973 11713 3007 11747
rect 3157 11713 3191 11747
rect 3709 11713 3743 11747
rect 3802 11713 3836 11747
rect 4077 11713 4111 11747
rect 4215 11713 4249 11747
rect 8033 11713 8067 11747
rect 8125 11713 8159 11747
rect 8309 11713 8343 11747
rect 8401 11713 8435 11747
rect 9309 11713 9343 11747
rect 9415 11713 9449 11747
rect 9781 11713 9815 11747
rect 9965 11713 9999 11747
rect 10147 11713 10181 11747
rect 12265 11713 12299 11747
rect 12449 11713 12483 11747
rect 12909 11713 12943 11747
rect 13093 11713 13127 11747
rect 14105 11713 14139 11747
rect 14289 11713 14323 11747
rect 14841 11713 14875 11747
rect 15025 11713 15059 11747
rect 16773 11713 16807 11747
rect 2697 11645 2731 11679
rect 2789 11645 2823 11679
rect 7113 11645 7147 11679
rect 7665 11577 7699 11611
rect 9321 11577 9355 11611
rect 12541 11577 12575 11611
rect 16957 11577 16991 11611
rect 6929 11509 6963 11543
rect 10333 11509 10367 11543
rect 14197 11509 14231 11543
rect 15117 11509 15151 11543
rect 3801 11305 3835 11339
rect 5273 11305 5307 11339
rect 6469 11305 6503 11339
rect 7573 11305 7607 11339
rect 8401 11305 8435 11339
rect 10425 11305 10459 11339
rect 11805 11305 11839 11339
rect 15209 11305 15243 11339
rect 17969 11305 18003 11339
rect 4169 11237 4203 11271
rect 6285 11237 6319 11271
rect 8217 11237 8251 11271
rect 8953 11237 8987 11271
rect 10241 11237 10275 11271
rect 11713 11237 11747 11271
rect 7757 11169 7791 11203
rect 7849 11169 7883 11203
rect 8493 11169 8527 11203
rect 12081 11169 12115 11203
rect 12265 11169 12299 11203
rect 15577 11169 15611 11203
rect 16221 11169 16255 11203
rect 1961 11101 1995 11135
rect 2145 11101 2179 11135
rect 2237 11101 2271 11135
rect 2605 11101 2639 11135
rect 2881 11101 2915 11135
rect 3985 11101 4019 11135
rect 4261 11101 4295 11135
rect 4997 11101 5031 11135
rect 5181 11101 5215 11135
rect 5457 11101 5491 11135
rect 5641 11101 5675 11135
rect 5917 11101 5951 11135
rect 6009 11101 6043 11135
rect 6285 11101 6319 11135
rect 6653 11101 6687 11135
rect 6745 11101 6779 11135
rect 6929 11101 6963 11135
rect 7021 11101 7055 11135
rect 7941 11101 7975 11135
rect 8033 11101 8067 11135
rect 8585 11101 8619 11135
rect 9229 11101 9263 11135
rect 9689 11101 9723 11135
rect 9873 11101 9907 11135
rect 10057 11101 10091 11135
rect 10149 11101 10183 11135
rect 11069 11101 11103 11135
rect 11162 11101 11196 11135
rect 11437 11101 11471 11135
rect 11534 11101 11568 11135
rect 11989 11101 12023 11135
rect 12173 11101 12207 11135
rect 13645 11101 13679 11135
rect 13829 11101 13863 11135
rect 13921 11101 13955 11135
rect 14105 11101 14139 11135
rect 14289 11101 14323 11135
rect 14381 11101 14415 11135
rect 14473 11101 14507 11135
rect 14749 11101 14783 11135
rect 15025 11101 15059 11135
rect 15301 11101 15335 11135
rect 15669 11101 15703 11135
rect 15853 11101 15887 11135
rect 3525 11033 3559 11067
rect 5089 11033 5123 11067
rect 5549 11033 5583 11067
rect 5779 11033 5813 11067
rect 6101 11033 6135 11067
rect 8953 11033 8987 11067
rect 9137 11033 9171 11067
rect 10609 11033 10643 11067
rect 11345 11033 11379 11067
rect 13461 11033 13495 11067
rect 14611 11033 14645 11067
rect 15393 11033 15427 11067
rect 15761 11033 15795 11067
rect 16497 11033 16531 11067
rect 2145 10965 2179 10999
rect 10409 10965 10443 10999
rect 14841 10965 14875 10999
rect 15485 10965 15519 10999
rect 16037 10965 16071 10999
rect 2605 10761 2639 10795
rect 5733 10761 5767 10795
rect 7021 10761 7055 10795
rect 9781 10761 9815 10795
rect 12449 10761 12483 10795
rect 12541 10761 12575 10795
rect 15301 10761 15335 10795
rect 16221 10761 16255 10795
rect 2881 10693 2915 10727
rect 2973 10693 3007 10727
rect 5365 10693 5399 10727
rect 12693 10693 12727 10727
rect 12909 10693 12943 10727
rect 16957 10693 16991 10727
rect 2789 10625 2823 10659
rect 3157 10625 3191 10659
rect 3249 10625 3283 10659
rect 3893 10625 3927 10659
rect 4537 10625 4571 10659
rect 4813 10625 4847 10659
rect 4997 10625 5031 10659
rect 5089 10625 5123 10659
rect 5182 10625 5216 10659
rect 5457 10625 5491 10659
rect 5595 10625 5629 10659
rect 6929 10625 6963 10659
rect 7113 10625 7147 10659
rect 8769 10625 8803 10659
rect 8953 10625 8987 10659
rect 9229 10625 9263 10659
rect 9321 10625 9355 10659
rect 9413 10625 9447 10659
rect 9960 10625 9994 10659
rect 10057 10625 10091 10659
rect 10149 10625 10183 10659
rect 10277 10625 10311 10659
rect 10425 10625 10459 10659
rect 10977 10625 11011 10659
rect 11161 10625 11195 10659
rect 11897 10625 11931 10659
rect 14013 10625 14047 10659
rect 14197 10625 14231 10659
rect 14289 10625 14323 10659
rect 14381 10625 14415 10659
rect 15485 10625 15519 10659
rect 15577 10625 15611 10659
rect 15761 10625 15795 10659
rect 15853 10625 15887 10659
rect 16313 10625 16347 10659
rect 17325 10625 17359 10659
rect 3985 10557 4019 10591
rect 4629 10557 4663 10591
rect 9137 10557 9171 10591
rect 12173 10557 12207 10591
rect 16840 10557 16874 10591
rect 17049 10557 17083 10591
rect 4721 10489 4755 10523
rect 11345 10489 11379 10523
rect 16681 10489 16715 10523
rect 3893 10421 3927 10455
rect 4261 10421 4295 10455
rect 4353 10421 4387 10455
rect 8861 10421 8895 10455
rect 9597 10421 9631 10455
rect 11069 10421 11103 10455
rect 12265 10421 12299 10455
rect 12725 10421 12759 10455
rect 14657 10421 14691 10455
rect 3341 10217 3375 10251
rect 6837 10217 6871 10251
rect 7481 10217 7515 10251
rect 9689 10217 9723 10251
rect 16221 10217 16255 10251
rect 16405 10217 16439 10251
rect 9229 10149 9263 10183
rect 16773 10149 16807 10183
rect 2697 10081 2731 10115
rect 2835 10081 2869 10115
rect 4077 10081 4111 10115
rect 4169 10081 4203 10115
rect 4261 10081 4295 10115
rect 6929 10081 6963 10115
rect 8677 10081 8711 10115
rect 9321 10081 9355 10115
rect 11161 10081 11195 10115
rect 11253 10081 11287 10115
rect 11621 10081 11655 10115
rect 2513 10013 2547 10047
rect 2973 10013 3007 10047
rect 3065 10013 3099 10047
rect 3341 10013 3375 10047
rect 3985 10013 4019 10047
rect 4629 10013 4663 10047
rect 4808 10013 4842 10047
rect 4905 10013 4939 10047
rect 4997 10013 5031 10047
rect 7021 10013 7055 10047
rect 7113 10013 7147 10047
rect 7297 10013 7331 10047
rect 8585 10013 8619 10047
rect 8769 10013 8803 10047
rect 8953 10013 8987 10047
rect 9137 10013 9171 10047
rect 9413 10013 9447 10047
rect 10885 10013 10919 10047
rect 11069 10013 11103 10047
rect 11437 10013 11471 10047
rect 11897 10013 11931 10047
rect 11989 10013 12023 10047
rect 12265 10013 12299 10047
rect 12357 10013 12391 10047
rect 12633 10013 12667 10047
rect 12817 10013 12851 10047
rect 13093 10013 13127 10047
rect 13460 10013 13494 10047
rect 13553 10013 13587 10047
rect 14656 10013 14690 10047
rect 14749 10013 14783 10047
rect 15393 10013 15427 10047
rect 15577 10013 15611 10047
rect 15945 10013 15979 10047
rect 16865 10013 16899 10047
rect 17233 10013 17267 10047
rect 3157 9945 3191 9979
rect 5733 9945 5767 9979
rect 6285 9945 6319 9979
rect 7573 9945 7607 9979
rect 9965 9945 9999 9979
rect 12081 9945 12115 9979
rect 12725 9945 12759 9979
rect 12955 9945 12989 9979
rect 14381 9945 14415 9979
rect 15301 9945 15335 9979
rect 16405 9945 16439 9979
rect 2513 9877 2547 9911
rect 3801 9877 3835 9911
rect 5273 9877 5307 9911
rect 5457 9877 5491 9911
rect 6009 9877 6043 9911
rect 6653 9877 6687 9911
rect 7297 9877 7331 9911
rect 9873 9877 9907 9911
rect 11713 9877 11747 9911
rect 12449 9877 12483 9911
rect 13185 9877 13219 9911
rect 16037 9877 16071 9911
rect 2973 9673 3007 9707
rect 3801 9673 3835 9707
rect 9873 9673 9907 9707
rect 14933 9673 14967 9707
rect 2329 9605 2363 9639
rect 4261 9605 4295 9639
rect 5457 9605 5491 9639
rect 5825 9605 5859 9639
rect 7849 9605 7883 9639
rect 12449 9605 12483 9639
rect 12541 9605 12575 9639
rect 16129 9605 16163 9639
rect 1685 9537 1719 9571
rect 2513 9537 2547 9571
rect 2605 9537 2639 9571
rect 2789 9537 2823 9571
rect 2881 9537 2915 9571
rect 3157 9537 3191 9571
rect 3249 9537 3283 9571
rect 3433 9537 3467 9571
rect 3525 9537 3559 9571
rect 3617 9537 3651 9571
rect 4445 9537 4479 9571
rect 4629 9537 4663 9571
rect 4721 9537 4755 9571
rect 5273 9537 5307 9571
rect 5641 9537 5675 9571
rect 5917 9537 5951 9571
rect 6561 9537 6595 9571
rect 6653 9537 6687 9571
rect 7297 9537 7331 9571
rect 7573 9537 7607 9571
rect 7757 9537 7791 9571
rect 9781 9537 9815 9571
rect 10149 9537 10183 9571
rect 12265 9537 12299 9571
rect 12633 9537 12667 9571
rect 13185 9537 13219 9571
rect 13913 9537 13947 9571
rect 14005 9537 14039 9571
rect 14197 9537 14231 9571
rect 14289 9537 14323 9571
rect 14381 9537 14415 9571
rect 14473 9537 14507 9571
rect 14657 9537 14691 9571
rect 14749 9537 14783 9571
rect 16681 9537 16715 9571
rect 17693 9537 17727 9571
rect 1777 9469 1811 9503
rect 2145 9469 2179 9503
rect 4905 9469 4939 9503
rect 4997 9469 5031 9503
rect 6745 9469 6779 9503
rect 6837 9469 6871 9503
rect 7205 9469 7239 9503
rect 7665 9469 7699 9503
rect 9965 9469 9999 9503
rect 16957 9469 16991 9503
rect 7021 9401 7055 9435
rect 13001 9401 13035 9435
rect 14657 9401 14691 9435
rect 1501 9333 1535 9367
rect 6377 9333 6411 9367
rect 10149 9333 10183 9367
rect 12817 9333 12851 9367
rect 13737 9333 13771 9367
rect 16405 9333 16439 9367
rect 17785 9333 17819 9367
rect 2329 9129 2363 9163
rect 2789 9129 2823 9163
rect 3271 9129 3305 9163
rect 6193 9129 6227 9163
rect 7757 9129 7791 9163
rect 9505 9129 9539 9163
rect 14381 9129 14415 9163
rect 3433 9061 3467 9095
rect 3801 9061 3835 9095
rect 4353 9061 4387 9095
rect 15025 9061 15059 9095
rect 6377 8993 6411 9027
rect 1685 8925 1719 8959
rect 2513 8925 2547 8959
rect 2605 8925 2639 8959
rect 4077 8925 4111 8959
rect 4169 8925 4203 8959
rect 4261 8925 4295 8959
rect 4537 8925 4571 8959
rect 6193 8925 6227 8959
rect 6469 8925 6503 8959
rect 6561 8925 6595 8959
rect 7573 8925 7607 8959
rect 8125 8925 8159 8959
rect 9229 8925 9263 8959
rect 9597 8925 9631 8959
rect 9781 8925 9815 8959
rect 9873 8925 9907 8959
rect 10057 8925 10091 8959
rect 10149 8925 10183 8959
rect 11805 8925 11839 8959
rect 12173 8925 12207 8959
rect 12265 8925 12299 8959
rect 14473 8925 14507 8959
rect 14749 8925 14783 8959
rect 14841 8925 14875 8959
rect 15209 8925 15243 8959
rect 15853 8925 15887 8959
rect 16129 8925 16163 8959
rect 16313 8925 16347 8959
rect 16589 8925 16623 8959
rect 17049 8925 17083 8959
rect 17417 8925 17451 8959
rect 2789 8857 2823 8891
rect 3065 8857 3099 8891
rect 4997 8857 5031 8891
rect 7941 8857 7975 8891
rect 9505 8857 9539 8891
rect 11897 8857 11931 8891
rect 11989 8857 12023 8891
rect 1501 8789 1535 8823
rect 3265 8789 3299 8823
rect 5089 8789 5123 8823
rect 7389 8789 7423 8823
rect 9321 8789 9355 8823
rect 11621 8789 11655 8823
rect 14197 8789 14231 8823
rect 15393 8789 15427 8823
rect 15669 8789 15703 8823
rect 15945 8789 15979 8823
rect 16681 8789 16715 8823
rect 4077 8585 4111 8619
rect 6377 8585 6411 8619
rect 14473 8585 14507 8619
rect 14933 8585 14967 8619
rect 16681 8585 16715 8619
rect 5825 8517 5859 8551
rect 6009 8517 6043 8551
rect 11529 8517 11563 8551
rect 12817 8517 12851 8551
rect 13185 8517 13219 8551
rect 4353 8449 4387 8483
rect 4445 8449 4479 8483
rect 5365 8449 5399 8483
rect 5549 8449 5583 8483
rect 6561 8449 6595 8483
rect 6745 8449 6779 8483
rect 7388 8449 7422 8483
rect 7665 8449 7699 8483
rect 7849 8449 7883 8483
rect 8125 8449 8159 8483
rect 8401 8449 8435 8483
rect 8585 8449 8619 8483
rect 8677 8449 8711 8483
rect 8861 8449 8895 8483
rect 9045 8449 9079 8483
rect 9229 8449 9263 8483
rect 9321 8449 9355 8483
rect 9413 8449 9447 8483
rect 10057 8449 10091 8483
rect 10149 8449 10183 8483
rect 10241 8449 10275 8483
rect 10425 8449 10459 8483
rect 10793 8449 10827 8483
rect 10885 8449 10919 8483
rect 11069 8449 11103 8483
rect 11161 8449 11195 8483
rect 11345 8449 11379 8483
rect 11785 8449 11819 8483
rect 11897 8449 11931 8483
rect 12010 8449 12044 8483
rect 12173 8449 12207 8483
rect 13001 8449 13035 8483
rect 13461 8449 13495 8483
rect 13737 8449 13771 8483
rect 14197 8449 14231 8483
rect 14289 8449 14323 8483
rect 14565 8449 14599 8483
rect 14749 8449 14783 8483
rect 14841 8449 14875 8483
rect 15117 8449 15151 8483
rect 15209 8449 15243 8483
rect 15301 8449 15335 8483
rect 15485 8449 15519 8483
rect 15577 8449 15611 8483
rect 15853 8449 15887 8483
rect 16129 8449 16163 8483
rect 16313 8449 16347 8483
rect 16497 8449 16531 8483
rect 16865 8449 16899 8483
rect 16957 8449 16991 8483
rect 5733 8381 5767 8415
rect 6653 8381 6687 8415
rect 6837 8381 6871 8415
rect 7113 8381 7147 8415
rect 7205 8381 7239 8415
rect 7297 8381 7331 8415
rect 13553 8381 13587 8415
rect 14013 8381 14047 8415
rect 14105 8381 14139 8415
rect 15669 8381 15703 8415
rect 16037 8381 16071 8415
rect 16405 8381 16439 8415
rect 6193 8313 6227 8347
rect 7573 8313 7607 8347
rect 7757 8313 7791 8347
rect 7941 8313 7975 8347
rect 8217 8313 8251 8347
rect 8309 8313 8343 8347
rect 8769 8313 8803 8347
rect 9689 8313 9723 8347
rect 9781 8313 9815 8347
rect 13645 8313 13679 8347
rect 15945 8313 15979 8347
rect 4445 8245 4479 8279
rect 13277 8245 13311 8279
rect 14565 8245 14599 8279
rect 2973 8041 3007 8075
rect 6469 8041 6503 8075
rect 7481 8041 7515 8075
rect 13369 8041 13403 8075
rect 14197 8041 14231 8075
rect 15945 8041 15979 8075
rect 2881 7973 2915 8007
rect 4537 7973 4571 8007
rect 4261 7905 4295 7939
rect 5089 7905 5123 7939
rect 6929 7905 6963 7939
rect 9137 7905 9171 7939
rect 11161 7905 11195 7939
rect 11621 7905 11655 7939
rect 11897 7905 11931 7939
rect 13277 7905 13311 7939
rect 13737 7905 13771 7939
rect 2789 7837 2823 7871
rect 3801 7837 3835 7871
rect 3985 7837 4019 7871
rect 4445 7837 4479 7871
rect 4629 7837 4663 7871
rect 5457 7837 5491 7871
rect 5549 7837 5583 7871
rect 5825 7837 5859 7871
rect 5973 7837 6007 7871
rect 6290 7837 6324 7871
rect 6745 7837 6779 7871
rect 7297 7837 7331 7871
rect 7389 7837 7423 7871
rect 7573 7837 7607 7871
rect 9229 7837 9263 7871
rect 9321 7837 9355 7871
rect 9413 7837 9447 7871
rect 9868 7837 9902 7871
rect 10057 7837 10091 7871
rect 10185 7837 10219 7871
rect 10333 7837 10367 7871
rect 11061 7837 11095 7871
rect 11253 7837 11287 7871
rect 11345 7837 11379 7871
rect 11529 7837 11563 7871
rect 11805 7837 11839 7871
rect 11989 7837 12023 7871
rect 12081 7837 12115 7871
rect 12265 7837 12299 7871
rect 13553 7837 13587 7871
rect 14105 7837 14139 7871
rect 14568 7837 14602 7871
rect 15761 7837 15795 7871
rect 15945 7837 15979 7871
rect 17785 7837 17819 7871
rect 3065 7769 3099 7803
rect 5733 7769 5767 7803
rect 6101 7769 6135 7803
rect 6193 7769 6227 7803
rect 9965 7769 9999 7803
rect 4077 7701 4111 7735
rect 6561 7701 6595 7735
rect 7113 7701 7147 7735
rect 9597 7701 9631 7735
rect 9689 7701 9723 7735
rect 10885 7701 10919 7735
rect 14565 7701 14599 7735
rect 14749 7701 14783 7735
rect 17969 7701 18003 7735
rect 3065 7497 3099 7531
rect 5825 7497 5859 7531
rect 10057 7497 10091 7531
rect 11989 7497 12023 7531
rect 15117 7497 15151 7531
rect 15853 7497 15887 7531
rect 2881 7429 2915 7463
rect 10885 7429 10919 7463
rect 2513 7361 2547 7395
rect 3525 7361 3559 7395
rect 3801 7361 3835 7395
rect 3985 7361 4019 7395
rect 4261 7361 4295 7395
rect 4353 7361 4387 7395
rect 4537 7361 4571 7395
rect 5641 7361 5675 7395
rect 7389 7361 7423 7395
rect 7665 7361 7699 7395
rect 7757 7361 7791 7395
rect 9229 7361 9263 7395
rect 9505 7361 9539 7395
rect 9689 7361 9723 7395
rect 10241 7361 10275 7395
rect 10333 7361 10367 7395
rect 10425 7361 10459 7395
rect 10563 7361 10597 7395
rect 10977 7361 11011 7395
rect 11805 7361 11839 7395
rect 12449 7361 12483 7395
rect 12633 7361 12667 7395
rect 12909 7361 12943 7395
rect 13001 7361 13035 7395
rect 13369 7361 13403 7395
rect 13553 7361 13587 7395
rect 13921 7361 13955 7395
rect 14105 7361 14139 7395
rect 15301 7361 15335 7395
rect 15577 7361 15611 7395
rect 15761 7361 15795 7395
rect 16221 7361 16255 7395
rect 17233 7361 17267 7395
rect 5365 7293 5399 7327
rect 5457 7293 5491 7327
rect 5549 7293 5583 7327
rect 7481 7293 7515 7327
rect 9045 7293 9079 7327
rect 9413 7293 9447 7327
rect 10701 7293 10735 7327
rect 11529 7293 11563 7327
rect 12817 7293 12851 7327
rect 13093 7293 13127 7327
rect 13277 7293 13311 7327
rect 13737 7293 13771 7327
rect 13829 7293 13863 7327
rect 15485 7293 15519 7327
rect 16129 7293 16163 7327
rect 17049 7293 17083 7327
rect 7941 7225 7975 7259
rect 9321 7225 9355 7259
rect 12541 7225 12575 7259
rect 15393 7225 15427 7259
rect 2881 7157 2915 7191
rect 3341 7157 3375 7191
rect 4077 7157 4111 7191
rect 4353 7157 4387 7191
rect 11621 7157 11655 7191
rect 16037 7157 16071 7191
rect 7021 6953 7055 6987
rect 6285 6885 6319 6919
rect 11897 6885 11931 6919
rect 16589 6885 16623 6919
rect 14197 6817 14231 6851
rect 14565 6817 14599 6851
rect 16405 6817 16439 6851
rect 5457 6749 5491 6783
rect 5549 6749 5583 6783
rect 5733 6749 5767 6783
rect 5825 6749 5859 6783
rect 7021 6749 7055 6783
rect 7297 6749 7331 6783
rect 7389 6749 7423 6783
rect 7573 6749 7607 6783
rect 7665 6749 7699 6783
rect 7849 6749 7883 6783
rect 11897 6749 11931 6783
rect 12081 6749 12115 6783
rect 14381 6749 14415 6783
rect 14473 6749 14507 6783
rect 14657 6749 14691 6783
rect 15117 6749 15151 6783
rect 15209 6749 15243 6783
rect 15301 6749 15335 6783
rect 15485 6749 15519 6783
rect 6009 6681 6043 6715
rect 7205 6681 7239 6715
rect 7481 6681 7515 6715
rect 16865 6681 16899 6715
rect 5273 6613 5307 6647
rect 7757 6613 7791 6647
rect 14841 6613 14875 6647
rect 7297 6409 7331 6443
rect 8861 6409 8895 6443
rect 12173 6409 12207 6443
rect 16037 6409 16071 6443
rect 17785 6409 17819 6443
rect 2881 6341 2915 6375
rect 3097 6341 3131 6375
rect 3341 6341 3375 6375
rect 3709 6341 3743 6375
rect 6929 6341 6963 6375
rect 9965 6341 9999 6375
rect 14381 6341 14415 6375
rect 14749 6341 14783 6375
rect 14933 6341 14967 6375
rect 15301 6341 15335 6375
rect 3525 6273 3559 6307
rect 3801 6273 3835 6307
rect 4169 6273 4203 6307
rect 4261 6273 4295 6307
rect 4905 6295 4939 6329
rect 5181 6273 5215 6307
rect 5365 6273 5399 6307
rect 5457 6273 5491 6307
rect 5549 6273 5583 6307
rect 6009 6273 6043 6307
rect 6193 6273 6227 6307
rect 6837 6273 6871 6307
rect 7113 6273 7147 6307
rect 7665 6273 7699 6307
rect 7941 6273 7975 6307
rect 8125 6273 8159 6307
rect 8309 6273 8343 6307
rect 8585 6273 8619 6307
rect 8769 6273 8803 6307
rect 9045 6273 9079 6307
rect 9137 6273 9171 6307
rect 9229 6273 9263 6307
rect 9413 6273 9447 6307
rect 9505 6273 9539 6307
rect 9873 6273 9907 6307
rect 10149 6273 10183 6307
rect 10609 6273 10643 6307
rect 10793 6273 10827 6307
rect 10885 6273 10919 6307
rect 11529 6273 11563 6307
rect 11713 6273 11747 6307
rect 11805 6273 11839 6307
rect 11897 6273 11931 6307
rect 12541 6273 12575 6307
rect 12633 6273 12667 6307
rect 12725 6273 12759 6307
rect 12909 6273 12943 6307
rect 13185 6273 13219 6307
rect 13277 6273 13311 6307
rect 13461 6273 13495 6307
rect 13553 6273 13587 6307
rect 14473 6273 14507 6307
rect 14565 6273 14599 6307
rect 14841 6273 14875 6307
rect 15117 6273 15151 6307
rect 15393 6273 15427 6307
rect 15853 6273 15887 6307
rect 16957 6273 16991 6307
rect 4077 6205 4111 6239
rect 4353 6205 4387 6239
rect 4813 6205 4847 6239
rect 7757 6205 7791 6239
rect 7849 6205 7883 6239
rect 8677 6205 8711 6239
rect 10333 6205 10367 6239
rect 17049 6205 17083 6239
rect 4537 6137 4571 6171
rect 7481 6137 7515 6171
rect 8217 6137 8251 6171
rect 10701 6137 10735 6171
rect 3065 6069 3099 6103
rect 3249 6069 3283 6103
rect 3893 6069 3927 6103
rect 4905 6069 4939 6103
rect 5825 6069 5859 6103
rect 6009 6069 6043 6103
rect 9689 6069 9723 6103
rect 11069 6069 11103 6103
rect 12265 6069 12299 6103
rect 13001 6069 13035 6103
rect 3433 5865 3467 5899
rect 4353 5865 4387 5899
rect 4813 5865 4847 5899
rect 9689 5865 9723 5899
rect 11253 5865 11287 5899
rect 12265 5865 12299 5899
rect 12541 5865 12575 5899
rect 13277 5865 13311 5899
rect 16957 5865 16991 5899
rect 8125 5797 8159 5831
rect 10517 5797 10551 5831
rect 14657 5797 14691 5831
rect 4445 5729 4479 5763
rect 5181 5729 5215 5763
rect 5825 5729 5859 5763
rect 7297 5729 7331 5763
rect 7665 5729 7699 5763
rect 8033 5729 8067 5763
rect 13185 5729 13219 5763
rect 15945 5729 15979 5763
rect 1685 5661 1719 5695
rect 3926 5661 3960 5695
rect 4997 5661 5031 5695
rect 5273 5661 5307 5695
rect 5457 5661 5491 5695
rect 5641 5661 5675 5695
rect 5733 5661 5767 5695
rect 5917 5661 5951 5695
rect 6101 5661 6135 5695
rect 6929 5661 6963 5695
rect 7113 5661 7147 5695
rect 7205 5661 7239 5695
rect 7481 5661 7515 5695
rect 7941 5661 7975 5695
rect 8217 5661 8251 5695
rect 8953 5661 8987 5695
rect 9137 5661 9171 5695
rect 9229 5661 9263 5695
rect 9321 5661 9355 5695
rect 9505 5661 9539 5695
rect 9873 5661 9907 5695
rect 9966 5661 10000 5695
rect 10149 5661 10183 5695
rect 10338 5661 10372 5695
rect 10609 5661 10643 5695
rect 10793 5661 10827 5695
rect 10885 5661 10919 5695
rect 10977 5661 11011 5695
rect 11713 5661 11747 5695
rect 11805 5661 11839 5695
rect 11989 5661 12023 5695
rect 12081 5661 12115 5695
rect 12449 5661 12483 5695
rect 12633 5661 12667 5695
rect 13648 5661 13682 5695
rect 14933 5661 14967 5695
rect 15117 5661 15151 5695
rect 15301 5661 15335 5695
rect 16037 5661 16071 5695
rect 16681 5661 16715 5695
rect 3249 5593 3283 5627
rect 7757 5593 7791 5627
rect 10241 5593 10275 5627
rect 14473 5593 14507 5627
rect 15209 5593 15243 5627
rect 16865 5593 16899 5627
rect 1501 5525 1535 5559
rect 3449 5525 3483 5559
rect 3617 5525 3651 5559
rect 3801 5525 3835 5559
rect 3985 5525 4019 5559
rect 13645 5525 13679 5559
rect 13829 5525 13863 5559
rect 15485 5525 15519 5559
rect 3985 5321 4019 5355
rect 8677 5321 8711 5355
rect 12173 5321 12207 5355
rect 13461 5321 13495 5355
rect 13987 5321 14021 5355
rect 14289 5321 14323 5355
rect 16405 5321 16439 5355
rect 13369 5253 13403 5287
rect 14197 5253 14231 5287
rect 4353 5185 4387 5219
rect 6745 5185 6779 5219
rect 6929 5185 6963 5219
rect 7021 5185 7055 5219
rect 7113 5185 7147 5219
rect 8861 5185 8895 5219
rect 9137 5185 9171 5219
rect 10333 5185 10367 5219
rect 10793 5185 10827 5219
rect 12449 5185 12483 5219
rect 12541 5185 12575 5219
rect 12725 5185 12759 5219
rect 13277 5185 13311 5219
rect 14289 5185 14323 5219
rect 14473 5185 14507 5219
rect 15209 5185 15243 5219
rect 15301 5185 15335 5219
rect 15393 5185 15427 5219
rect 15577 5185 15611 5219
rect 15853 5185 15887 5219
rect 15945 5185 15979 5219
rect 16129 5185 16163 5219
rect 16221 5185 16255 5219
rect 16497 5185 16531 5219
rect 4261 5117 4295 5151
rect 8769 5117 8803 5151
rect 10517 5117 10551 5151
rect 12173 5117 12207 5151
rect 13645 5117 13679 5151
rect 13737 5117 13771 5151
rect 15669 5117 15703 5151
rect 10425 5049 10459 5083
rect 12909 5049 12943 5083
rect 15025 5049 15059 5083
rect 4353 4981 4387 5015
rect 7389 4981 7423 5015
rect 9045 4981 9079 5015
rect 10057 4981 10091 5015
rect 10609 4981 10643 5015
rect 12357 4981 12391 5015
rect 12541 4981 12575 5015
rect 13001 4981 13035 5015
rect 13829 4981 13863 5015
rect 14013 4981 14047 5015
rect 5733 4777 5767 4811
rect 11345 4777 11379 4811
rect 11989 4777 12023 4811
rect 12173 4777 12207 4811
rect 15761 4777 15795 4811
rect 15945 4777 15979 4811
rect 3341 4709 3375 4743
rect 15209 4709 15243 4743
rect 15393 4709 15427 4743
rect 6561 4641 6595 4675
rect 7113 4641 7147 4675
rect 7665 4641 7699 4675
rect 11437 4641 11471 4675
rect 15669 4641 15703 4675
rect 5457 4573 5491 4607
rect 5641 4573 5675 4607
rect 5917 4573 5951 4607
rect 6009 4573 6043 4607
rect 6469 4573 6503 4607
rect 6837 4573 6871 4607
rect 6929 4573 6963 4607
rect 7205 4573 7239 4607
rect 7389 4573 7423 4607
rect 7481 4573 7515 4607
rect 7757 4573 7791 4607
rect 11529 4573 11563 4607
rect 13277 4573 13311 4607
rect 13461 4573 13495 4607
rect 13829 4573 13863 4607
rect 14381 4573 14415 4607
rect 16313 4573 16347 4607
rect 2973 4505 3007 4539
rect 5273 4505 5307 4539
rect 5733 4505 5767 4539
rect 11805 4505 11839 4539
rect 15945 4505 15979 4539
rect 3433 4437 3467 4471
rect 6745 4437 6779 4471
rect 7205 4437 7239 4471
rect 11161 4437 11195 4471
rect 12005 4437 12039 4471
rect 13369 4437 13403 4471
rect 13645 4437 13679 4471
rect 14197 4437 14231 4471
rect 5733 4233 5767 4267
rect 6469 4233 6503 4267
rect 8585 4233 8619 4267
rect 8953 4233 8987 4267
rect 10977 4233 11011 4267
rect 11989 4233 12023 4267
rect 13093 4233 13127 4267
rect 4721 4165 4755 4199
rect 6009 4165 6043 4199
rect 6653 4165 6687 4199
rect 8769 4165 8803 4199
rect 13369 4165 13403 4199
rect 15025 4165 15059 4199
rect 3157 4097 3191 4131
rect 3433 4097 3467 4131
rect 5365 4097 5399 4131
rect 5825 4097 5859 4131
rect 6193 4097 6227 4131
rect 6377 4097 6411 4131
rect 6929 4097 6963 4131
rect 7205 4097 7239 4131
rect 7389 4097 7423 4131
rect 7757 4097 7791 4131
rect 8217 4097 8251 4131
rect 8401 4097 8435 4131
rect 8677 4097 8711 4131
rect 9045 4097 9079 4131
rect 9137 4097 9171 4131
rect 9229 4097 9263 4131
rect 9321 4097 9355 4131
rect 9597 4097 9631 4131
rect 9781 4097 9815 4131
rect 9873 4097 9907 4131
rect 9965 4097 9999 4131
rect 10149 4097 10183 4131
rect 10609 4097 10643 4131
rect 10793 4097 10827 4131
rect 11069 4097 11103 4131
rect 11713 4097 11747 4131
rect 11897 4097 11931 4131
rect 11989 4097 12023 4131
rect 12173 4097 12207 4131
rect 13277 4097 13311 4131
rect 13461 4097 13495 4131
rect 13645 4097 13679 4131
rect 13737 4097 13771 4131
rect 14933 4097 14967 4131
rect 15669 4097 15703 4131
rect 15945 4097 15979 4131
rect 16773 4097 16807 4131
rect 16865 4097 16899 4131
rect 17049 4097 17083 4131
rect 5181 4029 5215 4063
rect 5457 4029 5491 4063
rect 7573 4029 7607 4063
rect 7849 4029 7883 4063
rect 7941 4029 7975 4063
rect 8033 4029 8067 4063
rect 11805 4029 11839 4063
rect 5089 3961 5123 3995
rect 6653 3961 6687 3995
rect 10057 3961 10091 3995
rect 16865 3961 16899 3995
rect 5549 3893 5583 3927
rect 6745 3893 6779 3927
rect 8769 3893 8803 3927
rect 9413 3893 9447 3927
rect 5641 3689 5675 3723
rect 8493 3689 8527 3723
rect 8585 3689 8619 3723
rect 9689 3689 9723 3723
rect 11989 3689 12023 3723
rect 14749 3689 14783 3723
rect 7481 3621 7515 3655
rect 9321 3621 9355 3655
rect 12173 3621 12207 3655
rect 12817 3621 12851 3655
rect 3065 3553 3099 3587
rect 4997 3553 5031 3587
rect 6101 3553 6135 3587
rect 8401 3553 8435 3587
rect 9413 3553 9447 3587
rect 10977 3553 11011 3587
rect 3433 3485 3467 3519
rect 3617 3485 3651 3519
rect 4077 3485 4111 3519
rect 4353 3485 4387 3519
rect 5365 3485 5399 3519
rect 5457 3485 5491 3519
rect 6561 3485 6595 3519
rect 6837 3485 6871 3519
rect 7297 3485 7331 3519
rect 7389 3485 7423 3519
rect 7941 3485 7975 3519
rect 8677 3485 8711 3519
rect 9229 3485 9263 3519
rect 9505 3485 9539 3519
rect 9873 3485 9907 3519
rect 9965 3485 9999 3519
rect 10149 3485 10183 3519
rect 10241 3485 10275 3519
rect 10609 3485 10643 3519
rect 10885 3485 10919 3519
rect 11161 3485 11195 3519
rect 11253 3485 11287 3519
rect 11529 3485 11563 3519
rect 11621 3485 11655 3519
rect 11805 3485 11839 3519
rect 12081 3485 12115 3519
rect 12357 3485 12391 3519
rect 12817 3485 12851 3519
rect 13001 3485 13035 3519
rect 13093 3485 13127 3519
rect 13185 3485 13219 3519
rect 13369 3485 13403 3519
rect 13737 3485 13771 3519
rect 14335 3485 14369 3519
rect 14473 3485 14507 3519
rect 14841 3485 14875 3519
rect 15209 3485 15243 3519
rect 15393 3485 15427 3519
rect 7113 3417 7147 3451
rect 10425 3417 10459 3451
rect 14105 3417 14139 3451
rect 15301 3417 15335 3451
rect 3157 3349 3191 3383
rect 4353 3349 4387 3383
rect 9045 3349 9079 3383
rect 10793 3349 10827 3383
rect 10977 3349 11011 3383
rect 12541 3349 12575 3383
rect 13369 3349 13403 3383
rect 7389 3145 7423 3179
rect 10425 3145 10459 3179
rect 10885 3145 10919 3179
rect 12265 3145 12299 3179
rect 6377 3077 6411 3111
rect 9689 3077 9723 3111
rect 12725 3077 12759 3111
rect 12909 3077 12943 3111
rect 13001 3077 13035 3111
rect 13277 3077 13311 3111
rect 7021 3009 7055 3043
rect 7114 3009 7148 3043
rect 9045 3009 9079 3043
rect 9229 3009 9263 3043
rect 9321 3009 9355 3043
rect 9413 3009 9447 3043
rect 9965 3009 9999 3043
rect 10149 3009 10183 3043
rect 10241 3009 10275 3043
rect 10333 3009 10367 3043
rect 10517 3009 10551 3043
rect 10701 3009 10735 3043
rect 10885 3009 10919 3043
rect 12173 3009 12207 3043
rect 12357 3009 12391 3043
rect 13113 3009 13147 3043
rect 13461 3009 13495 3043
rect 13553 3009 13587 3043
rect 9781 2941 9815 2975
rect 13277 2941 13311 2975
rect 6653 2873 6687 2907
rect 6837 2805 6871 2839
rect 12725 2805 12759 2839
rect 9597 2601 9631 2635
rect 6837 2397 6871 2431
rect 9137 2397 9171 2431
rect 9505 2397 9539 2431
rect 9689 2397 9723 2431
rect 9781 2397 9815 2431
rect 13645 2397 13679 2431
rect 6653 2261 6687 2295
rect 9321 2261 9355 2295
rect 9965 2261 9999 2295
rect 13829 2261 13863 2295
<< metal1 >>
rect 1104 19066 18400 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 18400 19066
rect 1104 18992 18400 19014
rect 8018 18912 8024 18964
rect 8076 18912 8082 18964
rect 8662 18912 8668 18964
rect 8720 18912 8726 18964
rect 9950 18912 9956 18964
rect 10008 18912 10014 18964
rect 10594 18912 10600 18964
rect 10652 18912 10658 18964
rect 10870 18912 10876 18964
rect 10928 18952 10934 18964
rect 11241 18955 11299 18961
rect 11241 18952 11253 18955
rect 10928 18924 11253 18952
rect 10928 18912 10934 18924
rect 11241 18921 11253 18924
rect 11287 18921 11299 18955
rect 11241 18915 11299 18921
rect 13170 18912 13176 18964
rect 13228 18952 13234 18964
rect 13817 18955 13875 18961
rect 13817 18952 13829 18955
rect 13228 18924 13829 18952
rect 13228 18912 13234 18924
rect 13817 18921 13829 18924
rect 13863 18921 13875 18955
rect 13817 18915 13875 18921
rect 7558 18708 7564 18760
rect 7616 18748 7622 18760
rect 7837 18751 7895 18757
rect 7837 18748 7849 18751
rect 7616 18720 7849 18748
rect 7616 18708 7622 18720
rect 7837 18717 7849 18720
rect 7883 18717 7895 18751
rect 7837 18711 7895 18717
rect 8478 18708 8484 18760
rect 8536 18708 8542 18760
rect 9122 18708 9128 18760
rect 9180 18748 9186 18760
rect 9769 18751 9827 18757
rect 9769 18748 9781 18751
rect 9180 18720 9781 18748
rect 9180 18708 9186 18720
rect 9769 18717 9781 18720
rect 9815 18717 9827 18751
rect 9769 18711 9827 18717
rect 10042 18708 10048 18760
rect 10100 18748 10106 18760
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 10100 18720 10425 18748
rect 10100 18708 10106 18720
rect 10413 18717 10425 18720
rect 10459 18717 10471 18751
rect 10413 18711 10471 18717
rect 11057 18751 11115 18757
rect 11057 18717 11069 18751
rect 11103 18748 11115 18751
rect 11238 18748 11244 18760
rect 11103 18720 11244 18748
rect 11103 18717 11115 18720
rect 11057 18711 11115 18717
rect 11238 18708 11244 18720
rect 11296 18708 11302 18760
rect 12342 18708 12348 18760
rect 12400 18748 12406 18760
rect 13633 18751 13691 18757
rect 13633 18748 13645 18751
rect 12400 18720 13645 18748
rect 12400 18708 12406 18720
rect 13633 18717 13645 18720
rect 13679 18717 13691 18751
rect 13633 18711 13691 18717
rect 14458 18708 14464 18760
rect 14516 18708 14522 18760
rect 13449 18683 13507 18689
rect 13449 18649 13461 18683
rect 13495 18680 13507 18683
rect 13495 18652 14688 18680
rect 13495 18649 13507 18652
rect 13449 18643 13507 18649
rect 9674 18572 9680 18624
rect 9732 18612 9738 18624
rect 13354 18612 13360 18624
rect 9732 18584 13360 18612
rect 9732 18572 9738 18584
rect 13354 18572 13360 18584
rect 13412 18572 13418 18624
rect 14660 18612 14688 18652
rect 14734 18640 14740 18692
rect 14792 18640 14798 18692
rect 16666 18680 16672 18692
rect 15962 18652 16672 18680
rect 16666 18640 16672 18652
rect 16724 18640 16730 18692
rect 16209 18615 16267 18621
rect 16209 18612 16221 18615
rect 14660 18584 16221 18612
rect 16209 18581 16221 18584
rect 16255 18581 16267 18615
rect 16209 18575 16267 18581
rect 1104 18522 18400 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 18400 18522
rect 1104 18448 18400 18470
rect 7558 18368 7564 18420
rect 7616 18368 7622 18420
rect 7944 18380 9536 18408
rect 7944 18284 7972 18380
rect 9508 18340 9536 18380
rect 10042 18368 10048 18420
rect 10100 18368 10106 18420
rect 11238 18368 11244 18420
rect 11296 18368 11302 18420
rect 12342 18368 12348 18420
rect 12400 18368 12406 18420
rect 13357 18411 13415 18417
rect 13357 18377 13369 18411
rect 13403 18377 13415 18411
rect 13357 18371 13415 18377
rect 10781 18343 10839 18349
rect 10781 18340 10793 18343
rect 9508 18312 10793 18340
rect 10781 18309 10793 18312
rect 10827 18340 10839 18343
rect 13372 18340 13400 18371
rect 14277 18343 14335 18349
rect 14277 18340 14289 18343
rect 10827 18312 12112 18340
rect 13372 18312 14289 18340
rect 10827 18309 10839 18312
rect 10781 18303 10839 18309
rect 7926 18232 7932 18284
rect 7984 18232 7990 18284
rect 8021 18275 8079 18281
rect 8021 18241 8033 18275
rect 8067 18272 8079 18275
rect 8389 18275 8447 18281
rect 8389 18272 8401 18275
rect 8067 18244 8401 18272
rect 8067 18241 8079 18244
rect 8021 18235 8079 18241
rect 8389 18241 8401 18244
rect 8435 18241 8447 18275
rect 8389 18235 8447 18241
rect 8573 18275 8631 18281
rect 8573 18241 8585 18275
rect 8619 18272 8631 18275
rect 8619 18244 8708 18272
rect 8619 18241 8631 18244
rect 8573 18235 8631 18241
rect 8110 18164 8116 18216
rect 8168 18164 8174 18216
rect 8680 18068 8708 18244
rect 8846 18232 8852 18284
rect 8904 18232 8910 18284
rect 8941 18275 8999 18281
rect 8941 18241 8953 18275
rect 8987 18241 8999 18275
rect 9125 18275 9183 18281
rect 9125 18272 9137 18275
rect 8941 18235 8999 18241
rect 9048 18244 9137 18272
rect 8754 18164 8760 18216
rect 8812 18204 8818 18216
rect 8956 18204 8984 18235
rect 8812 18176 8984 18204
rect 9048 18204 9076 18244
rect 9125 18241 9137 18244
rect 9171 18241 9183 18275
rect 9125 18235 9183 18241
rect 9214 18232 9220 18284
rect 9272 18272 9278 18284
rect 9272 18244 9352 18272
rect 9272 18232 9278 18244
rect 9048 18176 9260 18204
rect 8812 18164 8818 18176
rect 9122 18096 9128 18148
rect 9180 18096 9186 18148
rect 9232 18145 9260 18176
rect 9217 18139 9275 18145
rect 9217 18105 9229 18139
rect 9263 18105 9275 18139
rect 9324 18136 9352 18244
rect 9398 18232 9404 18284
rect 9456 18232 9462 18284
rect 9493 18275 9551 18281
rect 9493 18241 9505 18275
rect 9539 18272 9551 18275
rect 9766 18272 9772 18284
rect 9539 18244 9772 18272
rect 9539 18241 9551 18244
rect 9493 18235 9551 18241
rect 9766 18232 9772 18244
rect 9824 18272 9830 18284
rect 9861 18275 9919 18281
rect 9861 18272 9873 18275
rect 9824 18244 9873 18272
rect 9824 18232 9830 18244
rect 9861 18241 9873 18244
rect 9907 18241 9919 18275
rect 9861 18235 9919 18241
rect 10042 18232 10048 18284
rect 10100 18272 10106 18284
rect 10873 18275 10931 18281
rect 10100 18244 10824 18272
rect 10100 18232 10106 18244
rect 9674 18164 9680 18216
rect 9732 18164 9738 18216
rect 10686 18164 10692 18216
rect 10744 18164 10750 18216
rect 10796 18204 10824 18244
rect 10873 18241 10885 18275
rect 10919 18272 10931 18275
rect 11517 18275 11575 18281
rect 11517 18272 11529 18275
rect 10919 18244 11529 18272
rect 10919 18241 10931 18244
rect 10873 18235 10931 18241
rect 11517 18241 11529 18244
rect 11563 18241 11575 18275
rect 11517 18235 11575 18241
rect 11698 18232 11704 18284
rect 11756 18232 11762 18284
rect 12084 18281 12112 18312
rect 14277 18309 14289 18312
rect 14323 18309 14335 18343
rect 16482 18340 16488 18352
rect 15502 18312 16488 18340
rect 14277 18303 14335 18309
rect 16482 18300 16488 18312
rect 16540 18300 16546 18352
rect 12069 18275 12127 18281
rect 12069 18241 12081 18275
rect 12115 18241 12127 18275
rect 12069 18235 12127 18241
rect 12986 18232 12992 18284
rect 13044 18232 13050 18284
rect 13538 18232 13544 18284
rect 13596 18232 13602 18284
rect 13630 18232 13636 18284
rect 13688 18232 13694 18284
rect 16025 18275 16083 18281
rect 16025 18241 16037 18275
rect 16071 18272 16083 18275
rect 16574 18272 16580 18284
rect 16071 18244 16580 18272
rect 16071 18241 16083 18244
rect 16025 18235 16083 18241
rect 16574 18232 16580 18244
rect 16632 18232 16638 18284
rect 11790 18204 11796 18216
rect 10796 18176 11796 18204
rect 11790 18164 11796 18176
rect 11848 18204 11854 18216
rect 11977 18207 12035 18213
rect 11977 18204 11989 18207
rect 11848 18176 11989 18204
rect 11848 18164 11854 18176
rect 11977 18173 11989 18176
rect 12023 18173 12035 18207
rect 11977 18167 12035 18173
rect 12342 18164 12348 18216
rect 12400 18164 12406 18216
rect 13081 18207 13139 18213
rect 13081 18173 13093 18207
rect 13127 18173 13139 18207
rect 13081 18167 13139 18173
rect 14001 18207 14059 18213
rect 14001 18173 14013 18207
rect 14047 18173 14059 18207
rect 14001 18167 14059 18173
rect 11698 18136 11704 18148
rect 9324 18108 11704 18136
rect 9217 18099 9275 18105
rect 11698 18096 11704 18108
rect 11756 18096 11762 18148
rect 13096 18136 13124 18167
rect 13722 18136 13728 18148
rect 13096 18108 13728 18136
rect 13722 18096 13728 18108
rect 13780 18096 13786 18148
rect 9674 18068 9680 18080
rect 8680 18040 9680 18068
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 10870 18028 10876 18080
rect 10928 18068 10934 18080
rect 11885 18071 11943 18077
rect 11885 18068 11897 18071
rect 10928 18040 11897 18068
rect 10928 18028 10934 18040
rect 11885 18037 11897 18040
rect 11931 18037 11943 18071
rect 11885 18031 11943 18037
rect 12158 18028 12164 18080
rect 12216 18028 12222 18080
rect 13814 18028 13820 18080
rect 13872 18028 13878 18080
rect 14016 18068 14044 18167
rect 15749 18139 15807 18145
rect 15749 18105 15761 18139
rect 15795 18136 15807 18139
rect 16758 18136 16764 18148
rect 15795 18108 16764 18136
rect 15795 18105 15807 18108
rect 15749 18099 15807 18105
rect 16758 18096 16764 18108
rect 16816 18096 16822 18148
rect 14458 18068 14464 18080
rect 14016 18040 14464 18068
rect 14458 18028 14464 18040
rect 14516 18028 14522 18080
rect 15838 18028 15844 18080
rect 15896 18068 15902 18080
rect 15933 18071 15991 18077
rect 15933 18068 15945 18071
rect 15896 18040 15945 18068
rect 15896 18028 15902 18040
rect 15933 18037 15945 18040
rect 15979 18037 15991 18071
rect 15933 18031 15991 18037
rect 1104 17978 18400 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 18400 17978
rect 1104 17904 18400 17926
rect 8846 17824 8852 17876
rect 8904 17864 8910 17876
rect 9398 17864 9404 17876
rect 8904 17836 9404 17864
rect 8904 17824 8910 17836
rect 9398 17824 9404 17836
rect 9456 17824 9462 17876
rect 9677 17867 9735 17873
rect 9677 17833 9689 17867
rect 9723 17864 9735 17867
rect 9766 17864 9772 17876
rect 9723 17836 9772 17864
rect 9723 17833 9735 17836
rect 9677 17827 9735 17833
rect 9766 17824 9772 17836
rect 9824 17824 9830 17876
rect 10042 17824 10048 17876
rect 10100 17824 10106 17876
rect 10686 17824 10692 17876
rect 10744 17824 10750 17876
rect 11514 17824 11520 17876
rect 11572 17864 11578 17876
rect 11977 17867 12035 17873
rect 11977 17864 11989 17867
rect 11572 17836 11989 17864
rect 11572 17824 11578 17836
rect 11977 17833 11989 17836
rect 12023 17833 12035 17867
rect 11977 17827 12035 17833
rect 12342 17824 12348 17876
rect 12400 17824 12406 17876
rect 13449 17867 13507 17873
rect 13449 17833 13461 17867
rect 13495 17864 13507 17867
rect 14734 17864 14740 17876
rect 13495 17836 14740 17864
rect 13495 17833 13507 17836
rect 13449 17827 13507 17833
rect 14734 17824 14740 17836
rect 14792 17824 14798 17876
rect 16666 17824 16672 17876
rect 16724 17824 16730 17876
rect 5718 17756 5724 17808
rect 5776 17796 5782 17808
rect 8202 17796 8208 17808
rect 5776 17768 8208 17796
rect 5776 17756 5782 17768
rect 8202 17756 8208 17768
rect 8260 17796 8266 17808
rect 9858 17796 9864 17808
rect 8260 17768 9864 17796
rect 8260 17756 8266 17768
rect 9858 17756 9864 17768
rect 9916 17756 9922 17808
rect 11793 17799 11851 17805
rect 11793 17765 11805 17799
rect 11839 17796 11851 17799
rect 12158 17796 12164 17808
rect 11839 17768 12164 17796
rect 11839 17765 11851 17768
rect 11793 17759 11851 17765
rect 12158 17756 12164 17768
rect 12216 17756 12222 17808
rect 13538 17796 13544 17808
rect 13280 17768 13544 17796
rect 9953 17731 10011 17737
rect 9953 17697 9965 17731
rect 9999 17728 10011 17731
rect 10594 17728 10600 17740
rect 9999 17700 10600 17728
rect 9999 17697 10011 17700
rect 9953 17691 10011 17697
rect 10594 17688 10600 17700
rect 10652 17688 10658 17740
rect 11698 17688 11704 17740
rect 11756 17728 11762 17740
rect 13280 17737 13308 17768
rect 13538 17756 13544 17768
rect 13596 17796 13602 17808
rect 14182 17796 14188 17808
rect 13596 17768 14188 17796
rect 13596 17756 13602 17768
rect 14182 17756 14188 17768
rect 14240 17756 14246 17808
rect 12069 17731 12127 17737
rect 12069 17728 12081 17731
rect 11756 17700 12081 17728
rect 11756 17688 11762 17700
rect 12069 17697 12081 17700
rect 12115 17697 12127 17731
rect 12069 17691 12127 17697
rect 13265 17731 13323 17737
rect 13265 17697 13277 17731
rect 13311 17697 13323 17731
rect 13265 17691 13323 17697
rect 13354 17688 13360 17740
rect 13412 17688 13418 17740
rect 13814 17688 13820 17740
rect 13872 17728 13878 17740
rect 14737 17731 14795 17737
rect 14737 17728 14749 17731
rect 13872 17700 14749 17728
rect 13872 17688 13878 17700
rect 14737 17697 14749 17700
rect 14783 17697 14795 17731
rect 14737 17691 14795 17697
rect 2038 17620 2044 17672
rect 2096 17660 2102 17672
rect 2593 17663 2651 17669
rect 2593 17660 2605 17663
rect 2096 17632 2605 17660
rect 2096 17620 2102 17632
rect 2593 17629 2605 17632
rect 2639 17660 2651 17663
rect 8754 17660 8760 17672
rect 2639 17632 8760 17660
rect 2639 17629 2651 17632
rect 2593 17623 2651 17629
rect 8754 17620 8760 17632
rect 8812 17660 8818 17672
rect 9214 17660 9220 17672
rect 8812 17632 9220 17660
rect 8812 17620 8818 17632
rect 9214 17620 9220 17632
rect 9272 17620 9278 17672
rect 10045 17663 10103 17669
rect 10045 17629 10057 17663
rect 10091 17660 10103 17663
rect 10870 17660 10876 17672
rect 10091 17632 10876 17660
rect 10091 17629 10103 17632
rect 10045 17623 10103 17629
rect 7926 17592 7932 17604
rect 2700 17564 7932 17592
rect 2498 17484 2504 17536
rect 2556 17524 2562 17536
rect 2700 17533 2728 17564
rect 7926 17552 7932 17564
rect 7984 17552 7990 17604
rect 9766 17552 9772 17604
rect 9824 17592 9830 17604
rect 10060 17592 10088 17623
rect 10870 17620 10876 17632
rect 10928 17620 10934 17672
rect 11517 17663 11575 17669
rect 11517 17629 11529 17663
rect 11563 17660 11575 17663
rect 11606 17660 11612 17672
rect 11563 17632 11612 17660
rect 11563 17629 11575 17632
rect 11517 17623 11575 17629
rect 11606 17620 11612 17632
rect 11664 17620 11670 17672
rect 11793 17663 11851 17669
rect 11793 17629 11805 17663
rect 11839 17660 11851 17663
rect 11974 17660 11980 17672
rect 11839 17632 11980 17660
rect 11839 17629 11851 17632
rect 11793 17623 11851 17629
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 13173 17663 13231 17669
rect 13173 17629 13185 17663
rect 13219 17660 13231 17663
rect 13372 17660 13400 17688
rect 13219 17632 13768 17660
rect 13219 17629 13231 17632
rect 13173 17623 13231 17629
rect 9824 17564 10088 17592
rect 10321 17595 10379 17601
rect 9824 17552 9830 17564
rect 10321 17561 10333 17595
rect 10367 17592 10379 17595
rect 10410 17592 10416 17604
rect 10367 17564 10416 17592
rect 10367 17561 10379 17564
rect 10321 17555 10379 17561
rect 10410 17552 10416 17564
rect 10468 17552 10474 17604
rect 10502 17552 10508 17604
rect 10560 17552 10566 17604
rect 12986 17592 12992 17604
rect 11440 17564 12992 17592
rect 2685 17527 2743 17533
rect 2685 17524 2697 17527
rect 2556 17496 2697 17524
rect 2556 17484 2562 17496
rect 2685 17493 2697 17496
rect 2731 17493 2743 17527
rect 2685 17487 2743 17493
rect 5994 17484 6000 17536
rect 6052 17524 6058 17536
rect 8018 17524 8024 17536
rect 6052 17496 8024 17524
rect 6052 17484 6058 17496
rect 8018 17484 8024 17496
rect 8076 17524 8082 17536
rect 11440 17524 11468 17564
rect 12986 17552 12992 17564
rect 13044 17592 13050 17604
rect 13354 17592 13360 17604
rect 13044 17564 13360 17592
rect 13044 17552 13050 17564
rect 13354 17552 13360 17564
rect 13412 17552 13418 17604
rect 13740 17592 13768 17632
rect 14458 17620 14464 17672
rect 14516 17620 14522 17672
rect 15838 17620 15844 17672
rect 15896 17620 15902 17672
rect 16574 17620 16580 17672
rect 16632 17660 16638 17672
rect 16761 17663 16819 17669
rect 16761 17660 16773 17663
rect 16632 17632 16773 17660
rect 16632 17620 16638 17632
rect 16761 17629 16773 17632
rect 16807 17629 16819 17663
rect 16761 17623 16819 17629
rect 13740 17564 14964 17592
rect 14936 17536 14964 17564
rect 16022 17552 16028 17604
rect 16080 17592 16086 17604
rect 16485 17595 16543 17601
rect 16485 17592 16497 17595
rect 16080 17564 16497 17592
rect 16080 17552 16086 17564
rect 16485 17561 16497 17564
rect 16531 17561 16543 17595
rect 16485 17555 16543 17561
rect 8076 17496 11468 17524
rect 8076 17484 8082 17496
rect 11514 17484 11520 17536
rect 11572 17524 11578 17536
rect 11609 17527 11667 17533
rect 11609 17524 11621 17527
rect 11572 17496 11621 17524
rect 11572 17484 11578 17496
rect 11609 17493 11621 17496
rect 11655 17493 11667 17527
rect 11609 17487 11667 17493
rect 14918 17484 14924 17536
rect 14976 17484 14982 17536
rect 1104 17434 18400 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 18400 17434
rect 1104 17360 18400 17382
rect 5718 17280 5724 17332
rect 5776 17280 5782 17332
rect 7009 17323 7067 17329
rect 7009 17289 7021 17323
rect 7055 17320 7067 17323
rect 7190 17320 7196 17332
rect 7055 17292 7196 17320
rect 7055 17289 7067 17292
rect 7009 17283 7067 17289
rect 7190 17280 7196 17292
rect 7248 17320 7254 17332
rect 7248 17292 8708 17320
rect 7248 17280 7254 17292
rect 4798 17252 4804 17264
rect 3896 17224 4804 17252
rect 3896 17193 3924 17224
rect 4798 17212 4804 17224
rect 4856 17212 4862 17264
rect 5828 17224 6868 17252
rect 5828 17196 5856 17224
rect 3881 17187 3939 17193
rect 3881 17153 3893 17187
rect 3927 17153 3939 17187
rect 3881 17147 3939 17153
rect 3973 17187 4031 17193
rect 3973 17153 3985 17187
rect 4019 17153 4031 17187
rect 3973 17147 4031 17153
rect 3418 17076 3424 17128
rect 3476 17116 3482 17128
rect 3988 17116 4016 17147
rect 4062 17144 4068 17196
rect 4120 17184 4126 17196
rect 5353 17187 5411 17193
rect 5353 17184 5365 17187
rect 4120 17156 5365 17184
rect 4120 17144 4126 17156
rect 5353 17153 5365 17156
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 3476 17088 4016 17116
rect 4157 17119 4215 17125
rect 3476 17076 3482 17088
rect 4157 17085 4169 17119
rect 4203 17116 4215 17119
rect 4614 17116 4620 17128
rect 4203 17088 4620 17116
rect 4203 17085 4215 17088
rect 4157 17079 4215 17085
rect 4614 17076 4620 17088
rect 4672 17076 4678 17128
rect 5368 17116 5396 17147
rect 5810 17144 5816 17196
rect 5868 17144 5874 17196
rect 5905 17187 5963 17193
rect 5905 17153 5917 17187
rect 5951 17184 5963 17187
rect 5994 17184 6000 17196
rect 5951 17156 6000 17184
rect 5951 17153 5963 17156
rect 5905 17147 5963 17153
rect 5920 17116 5948 17147
rect 5994 17144 6000 17156
rect 6052 17144 6058 17196
rect 6840 17193 6868 17224
rect 7300 17224 8524 17252
rect 7300 17193 7328 17224
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 6825 17187 6883 17193
rect 6825 17153 6837 17187
rect 6871 17184 6883 17187
rect 7285 17187 7343 17193
rect 7285 17184 7297 17187
rect 6871 17156 7297 17184
rect 6871 17153 6883 17156
rect 6825 17147 6883 17153
rect 7285 17153 7297 17156
rect 7331 17153 7343 17187
rect 7285 17147 7343 17153
rect 5368 17088 5948 17116
rect 5534 17008 5540 17060
rect 5592 17048 5598 17060
rect 5997 17051 6055 17057
rect 5997 17048 6009 17051
rect 5592 17020 6009 17048
rect 5592 17008 5598 17020
rect 5997 17017 6009 17020
rect 6043 17048 6055 17051
rect 6564 17048 6592 17147
rect 8018 17144 8024 17196
rect 8076 17144 8082 17196
rect 7466 17076 7472 17128
rect 7524 17116 7530 17128
rect 7653 17119 7711 17125
rect 7653 17116 7665 17119
rect 7524 17088 7665 17116
rect 7524 17076 7530 17088
rect 7653 17085 7665 17088
rect 7699 17085 7711 17119
rect 8496 17116 8524 17224
rect 8570 17144 8576 17196
rect 8628 17144 8634 17196
rect 8680 17193 8708 17292
rect 10410 17280 10416 17332
rect 10468 17280 10474 17332
rect 10870 17280 10876 17332
rect 10928 17280 10934 17332
rect 11790 17280 11796 17332
rect 11848 17320 11854 17332
rect 12434 17320 12440 17332
rect 11848 17292 12440 17320
rect 11848 17280 11854 17292
rect 12434 17280 12440 17292
rect 12492 17280 12498 17332
rect 13630 17280 13636 17332
rect 13688 17320 13694 17332
rect 13725 17323 13783 17329
rect 13725 17320 13737 17323
rect 13688 17292 13737 17320
rect 13688 17280 13694 17292
rect 13725 17289 13737 17292
rect 13771 17289 13783 17323
rect 13725 17283 13783 17289
rect 14182 17280 14188 17332
rect 14240 17280 14246 17332
rect 8846 17212 8852 17264
rect 8904 17252 8910 17264
rect 9033 17255 9091 17261
rect 9033 17252 9045 17255
rect 8904 17224 9045 17252
rect 8904 17212 8910 17224
rect 9033 17221 9045 17224
rect 9079 17221 9091 17255
rect 10045 17255 10103 17261
rect 10045 17252 10057 17255
rect 9033 17215 9091 17221
rect 9232 17224 10057 17252
rect 8665 17187 8723 17193
rect 8665 17153 8677 17187
rect 8711 17153 8723 17187
rect 8665 17147 8723 17153
rect 8938 17144 8944 17196
rect 8996 17184 9002 17196
rect 9232 17184 9260 17224
rect 10045 17221 10057 17224
rect 10091 17221 10103 17255
rect 10045 17215 10103 17221
rect 10318 17212 10324 17264
rect 10376 17252 10382 17264
rect 11057 17255 11115 17261
rect 11057 17252 11069 17255
rect 10376 17224 11069 17252
rect 10376 17212 10382 17224
rect 11057 17221 11069 17224
rect 11103 17252 11115 17255
rect 11103 17224 13492 17252
rect 11103 17221 11115 17224
rect 11057 17215 11115 17221
rect 8996 17156 9260 17184
rect 9493 17187 9551 17193
rect 8996 17144 9002 17156
rect 9493 17153 9505 17187
rect 9539 17184 9551 17187
rect 9858 17184 9864 17196
rect 9539 17156 9864 17184
rect 9539 17153 9551 17156
rect 9493 17147 9551 17153
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 10134 17144 10140 17196
rect 10192 17144 10198 17196
rect 10229 17187 10287 17193
rect 10229 17153 10241 17187
rect 10275 17153 10287 17187
rect 10229 17147 10287 17153
rect 8496 17088 9168 17116
rect 7653 17079 7711 17085
rect 9030 17048 9036 17060
rect 6043 17020 9036 17048
rect 6043 17017 6055 17020
rect 5997 17011 6055 17017
rect 9030 17008 9036 17020
rect 9088 17008 9094 17060
rect 3786 16940 3792 16992
rect 3844 16980 3850 16992
rect 7006 16980 7012 16992
rect 3844 16952 7012 16980
rect 3844 16940 3850 16952
rect 7006 16940 7012 16952
rect 7064 16940 7070 16992
rect 8389 16983 8447 16989
rect 8389 16949 8401 16983
rect 8435 16980 8447 16983
rect 8846 16980 8852 16992
rect 8435 16952 8852 16980
rect 8435 16949 8447 16952
rect 8389 16943 8447 16949
rect 8846 16940 8852 16952
rect 8904 16940 8910 16992
rect 9140 16980 9168 17088
rect 9214 17076 9220 17128
rect 9272 17076 9278 17128
rect 9766 17076 9772 17128
rect 9824 17076 9830 17128
rect 10244 17116 10272 17147
rect 10594 17144 10600 17196
rect 10652 17144 10658 17196
rect 11241 17187 11299 17193
rect 11241 17153 11253 17187
rect 11287 17184 11299 17187
rect 11606 17184 11612 17196
rect 11287 17156 11612 17184
rect 11287 17153 11299 17156
rect 11241 17147 11299 17153
rect 11606 17144 11612 17156
rect 11664 17144 11670 17196
rect 11790 17144 11796 17196
rect 11848 17144 11854 17196
rect 12250 17144 12256 17196
rect 12308 17184 12314 17196
rect 12308 17156 13308 17184
rect 12308 17144 12314 17156
rect 11054 17116 11060 17128
rect 10244 17088 11060 17116
rect 11054 17076 11060 17088
rect 11112 17076 11118 17128
rect 13280 17125 13308 17156
rect 13354 17144 13360 17196
rect 13412 17144 13418 17196
rect 13464 17128 13492 17224
rect 16758 17212 16764 17264
rect 16816 17212 16822 17264
rect 13722 17144 13728 17196
rect 13780 17184 13786 17196
rect 13817 17187 13875 17193
rect 13817 17184 13829 17187
rect 13780 17156 13829 17184
rect 13780 17144 13786 17156
rect 13817 17153 13829 17156
rect 13863 17153 13875 17187
rect 13817 17147 13875 17153
rect 14001 17187 14059 17193
rect 14001 17153 14013 17187
rect 14047 17184 14059 17187
rect 15102 17184 15108 17196
rect 14047 17156 15108 17184
rect 14047 17153 14059 17156
rect 14001 17147 14059 17153
rect 15102 17144 15108 17156
rect 15160 17144 15166 17196
rect 15194 17144 15200 17196
rect 15252 17184 15258 17196
rect 16485 17187 16543 17193
rect 16485 17184 16497 17187
rect 15252 17156 16497 17184
rect 15252 17144 15258 17156
rect 16485 17153 16497 17156
rect 16531 17153 16543 17187
rect 16485 17147 16543 17153
rect 11517 17119 11575 17125
rect 11517 17085 11529 17119
rect 11563 17085 11575 17119
rect 11517 17079 11575 17085
rect 13265 17119 13323 17125
rect 13265 17085 13277 17119
rect 13311 17085 13323 17119
rect 13265 17079 13323 17085
rect 9232 17048 9260 17076
rect 11422 17048 11428 17060
rect 9232 17020 11428 17048
rect 11422 17008 11428 17020
rect 11480 17048 11486 17060
rect 11532 17048 11560 17079
rect 11480 17020 11560 17048
rect 11480 17008 11486 17020
rect 11790 17008 11796 17060
rect 11848 17048 11854 17060
rect 13170 17048 13176 17060
rect 11848 17020 13176 17048
rect 11848 17008 11854 17020
rect 13170 17008 13176 17020
rect 13228 17008 13234 17060
rect 13280 17048 13308 17079
rect 13446 17076 13452 17128
rect 13504 17076 13510 17128
rect 13541 17119 13599 17125
rect 13541 17085 13553 17119
rect 13587 17116 13599 17119
rect 13630 17116 13636 17128
rect 13587 17088 13636 17116
rect 13587 17085 13599 17088
rect 13541 17079 13599 17085
rect 13630 17076 13636 17088
rect 13688 17076 13694 17128
rect 14090 17076 14096 17128
rect 14148 17116 14154 17128
rect 14458 17116 14464 17128
rect 14148 17088 14464 17116
rect 14148 17076 14154 17088
rect 14458 17076 14464 17088
rect 14516 17116 14522 17128
rect 14737 17119 14795 17125
rect 14737 17116 14749 17119
rect 14516 17088 14749 17116
rect 14516 17076 14522 17088
rect 14737 17085 14749 17088
rect 14783 17085 14795 17119
rect 14737 17079 14795 17085
rect 14642 17048 14648 17060
rect 13280 17020 14648 17048
rect 14642 17008 14648 17020
rect 14700 17048 14706 17060
rect 16022 17048 16028 17060
rect 14700 17020 16028 17048
rect 14700 17008 14706 17020
rect 16022 17008 16028 17020
rect 16080 17008 16086 17060
rect 10410 16980 10416 16992
rect 9140 16952 10416 16980
rect 10410 16940 10416 16952
rect 10468 16980 10474 16992
rect 10689 16983 10747 16989
rect 10689 16980 10701 16983
rect 10468 16952 10701 16980
rect 10468 16940 10474 16952
rect 10689 16949 10701 16952
rect 10735 16949 10747 16983
rect 10689 16943 10747 16949
rect 13354 16940 13360 16992
rect 13412 16980 13418 16992
rect 16206 16980 16212 16992
rect 13412 16952 16212 16980
rect 13412 16940 13418 16952
rect 16206 16940 16212 16952
rect 16264 16980 16270 16992
rect 16853 16983 16911 16989
rect 16853 16980 16865 16983
rect 16264 16952 16865 16980
rect 16264 16940 16270 16952
rect 16853 16949 16865 16952
rect 16899 16949 16911 16983
rect 16853 16943 16911 16949
rect 1104 16890 18400 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 18400 16890
rect 1104 16816 18400 16838
rect 7653 16779 7711 16785
rect 7653 16745 7665 16779
rect 7699 16776 7711 16779
rect 8110 16776 8116 16788
rect 7699 16748 8116 16776
rect 7699 16745 7711 16748
rect 7653 16739 7711 16745
rect 8110 16736 8116 16748
rect 8168 16736 8174 16788
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 10321 16779 10379 16785
rect 10321 16776 10333 16779
rect 9916 16748 10333 16776
rect 9916 16736 9922 16748
rect 10321 16745 10333 16748
rect 10367 16745 10379 16779
rect 10321 16739 10379 16745
rect 13722 16736 13728 16788
rect 13780 16736 13786 16788
rect 15102 16736 15108 16788
rect 15160 16736 15166 16788
rect 5169 16711 5227 16717
rect 5169 16708 5181 16711
rect 3988 16680 5181 16708
rect 3605 16643 3663 16649
rect 3605 16609 3617 16643
rect 3651 16640 3663 16643
rect 3786 16640 3792 16652
rect 3651 16612 3792 16640
rect 3651 16609 3663 16612
rect 3605 16603 3663 16609
rect 3786 16600 3792 16612
rect 3844 16600 3850 16652
rect 3988 16649 4016 16680
rect 5169 16677 5181 16680
rect 5215 16677 5227 16711
rect 5626 16708 5632 16720
rect 5169 16671 5227 16677
rect 5276 16680 5632 16708
rect 3973 16643 4031 16649
rect 3973 16609 3985 16643
rect 4019 16609 4031 16643
rect 3973 16603 4031 16609
rect 4062 16600 4068 16652
rect 4120 16600 4126 16652
rect 4157 16643 4215 16649
rect 4157 16609 4169 16643
rect 4203 16640 4215 16643
rect 4525 16643 4583 16649
rect 4525 16640 4537 16643
rect 4203 16612 4537 16640
rect 4203 16609 4215 16612
rect 4157 16603 4215 16609
rect 4525 16609 4537 16612
rect 4571 16609 4583 16643
rect 5276 16640 5304 16680
rect 5626 16668 5632 16680
rect 5684 16668 5690 16720
rect 7006 16668 7012 16720
rect 7064 16708 7070 16720
rect 7064 16680 7972 16708
rect 7064 16668 7070 16680
rect 4525 16603 4583 16609
rect 4632 16612 5304 16640
rect 2590 16532 2596 16584
rect 2648 16572 2654 16584
rect 3237 16575 3295 16581
rect 3237 16572 3249 16575
rect 2648 16544 3249 16572
rect 2648 16532 2654 16544
rect 3237 16541 3249 16544
rect 3283 16541 3295 16575
rect 3237 16535 3295 16541
rect 3418 16532 3424 16584
rect 3476 16532 3482 16584
rect 4249 16575 4307 16581
rect 4249 16541 4261 16575
rect 4295 16572 4307 16575
rect 4632 16572 4660 16612
rect 5350 16600 5356 16652
rect 5408 16600 5414 16652
rect 5534 16600 5540 16652
rect 5592 16600 5598 16652
rect 7944 16649 7972 16680
rect 8570 16668 8576 16720
rect 8628 16708 8634 16720
rect 11790 16708 11796 16720
rect 8628 16680 11796 16708
rect 8628 16668 8634 16680
rect 11790 16668 11796 16680
rect 11848 16668 11854 16720
rect 13081 16711 13139 16717
rect 13081 16677 13093 16711
rect 13127 16708 13139 16711
rect 15010 16708 15016 16720
rect 13127 16680 15016 16708
rect 13127 16677 13139 16680
rect 13081 16671 13139 16677
rect 15010 16668 15016 16680
rect 15068 16668 15074 16720
rect 7193 16643 7251 16649
rect 7193 16609 7205 16643
rect 7239 16640 7251 16643
rect 7745 16643 7803 16649
rect 7745 16640 7757 16643
rect 7239 16612 7757 16640
rect 7239 16609 7251 16612
rect 7193 16603 7251 16609
rect 7745 16609 7757 16612
rect 7791 16609 7803 16643
rect 7745 16603 7803 16609
rect 7929 16643 7987 16649
rect 7929 16609 7941 16643
rect 7975 16609 7987 16643
rect 7929 16603 7987 16609
rect 8021 16643 8079 16649
rect 8021 16609 8033 16643
rect 8067 16609 8079 16643
rect 8021 16603 8079 16609
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16640 8263 16643
rect 9582 16640 9588 16652
rect 8251 16612 9588 16640
rect 8251 16609 8263 16612
rect 8205 16603 8263 16609
rect 4295 16544 4660 16572
rect 4295 16541 4307 16544
rect 4249 16535 4307 16541
rect 4706 16532 4712 16584
rect 4764 16532 4770 16584
rect 4798 16532 4804 16584
rect 4856 16532 4862 16584
rect 4982 16532 4988 16584
rect 5040 16532 5046 16584
rect 5077 16575 5135 16581
rect 5077 16541 5089 16575
rect 5123 16572 5135 16575
rect 5258 16572 5264 16584
rect 5123 16544 5264 16572
rect 5123 16541 5135 16544
rect 5077 16535 5135 16541
rect 5258 16532 5264 16544
rect 5316 16572 5322 16584
rect 5445 16575 5503 16581
rect 5445 16572 5457 16575
rect 5316 16544 5457 16572
rect 5316 16532 5322 16544
rect 5445 16541 5457 16544
rect 5491 16541 5503 16575
rect 5445 16535 5503 16541
rect 5629 16575 5687 16581
rect 5629 16541 5641 16575
rect 5675 16572 5687 16575
rect 5902 16572 5908 16584
rect 5675 16544 5908 16572
rect 5675 16541 5687 16544
rect 5629 16535 5687 16541
rect 5902 16532 5908 16544
rect 5960 16532 5966 16584
rect 6086 16532 6092 16584
rect 6144 16532 6150 16584
rect 6917 16575 6975 16581
rect 6917 16572 6929 16575
rect 6196 16544 6929 16572
rect 3050 16464 3056 16516
rect 3108 16504 3114 16516
rect 3436 16504 3464 16532
rect 6196 16504 6224 16544
rect 6917 16541 6929 16544
rect 6963 16541 6975 16575
rect 6917 16535 6975 16541
rect 7098 16532 7104 16584
rect 7156 16532 7162 16584
rect 7285 16575 7343 16581
rect 7285 16541 7297 16575
rect 7331 16572 7343 16575
rect 7374 16572 7380 16584
rect 7331 16544 7380 16572
rect 7331 16541 7343 16544
rect 7285 16535 7343 16541
rect 7374 16532 7380 16544
rect 7432 16532 7438 16584
rect 7466 16532 7472 16584
rect 7524 16532 7530 16584
rect 3108 16476 3464 16504
rect 4448 16476 6224 16504
rect 3108 16464 3114 16476
rect 4448 16445 4476 16476
rect 6454 16464 6460 16516
rect 6512 16464 6518 16516
rect 6546 16464 6552 16516
rect 6604 16504 6610 16516
rect 6641 16507 6699 16513
rect 6641 16504 6653 16507
rect 6604 16476 6653 16504
rect 6604 16464 6610 16476
rect 6641 16473 6653 16476
rect 6687 16473 6699 16507
rect 8036 16504 8064 16603
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 10137 16643 10195 16649
rect 10137 16640 10149 16643
rect 9690 16612 10149 16640
rect 8110 16532 8116 16584
rect 8168 16532 8174 16584
rect 8754 16532 8760 16584
rect 8812 16532 8818 16584
rect 8941 16575 8999 16581
rect 8941 16541 8953 16575
rect 8987 16541 8999 16575
rect 8941 16535 8999 16541
rect 8956 16504 8984 16535
rect 9306 16532 9312 16584
rect 9364 16572 9370 16584
rect 9690 16572 9718 16612
rect 10137 16609 10149 16612
rect 10183 16609 10195 16643
rect 10137 16603 10195 16609
rect 10594 16600 10600 16652
rect 10652 16640 10658 16652
rect 12250 16640 12256 16652
rect 10652 16612 12256 16640
rect 10652 16600 10658 16612
rect 9364 16544 9718 16572
rect 9364 16532 9370 16544
rect 9766 16532 9772 16584
rect 9824 16572 9830 16584
rect 9861 16575 9919 16581
rect 9861 16572 9873 16575
rect 9824 16544 9873 16572
rect 9824 16532 9830 16544
rect 9861 16541 9873 16544
rect 9907 16541 9919 16575
rect 9861 16535 9919 16541
rect 9950 16532 9956 16584
rect 10008 16572 10014 16584
rect 10229 16575 10287 16581
rect 10229 16572 10241 16575
rect 10008 16544 10241 16572
rect 10008 16532 10014 16544
rect 10229 16541 10241 16544
rect 10275 16572 10287 16575
rect 10318 16572 10324 16584
rect 10275 16544 10324 16572
rect 10275 16541 10287 16544
rect 10229 16535 10287 16541
rect 10318 16532 10324 16544
rect 10376 16532 10382 16584
rect 10413 16575 10471 16581
rect 10413 16541 10425 16575
rect 10459 16572 10471 16575
rect 10502 16572 10508 16584
rect 10459 16544 10508 16572
rect 10459 16541 10471 16544
rect 10413 16535 10471 16541
rect 10502 16532 10508 16544
rect 10560 16532 10566 16584
rect 10796 16581 10824 16612
rect 12250 16600 12256 16612
rect 12308 16600 12314 16652
rect 13906 16640 13912 16652
rect 13556 16612 13912 16640
rect 10781 16575 10839 16581
rect 10781 16541 10793 16575
rect 10827 16541 10839 16575
rect 10781 16535 10839 16541
rect 11057 16575 11115 16581
rect 11057 16541 11069 16575
rect 11103 16572 11115 16575
rect 11238 16572 11244 16584
rect 11103 16544 11244 16572
rect 11103 16541 11115 16544
rect 11057 16535 11115 16541
rect 6641 16467 6699 16473
rect 6748 16476 8984 16504
rect 4433 16439 4491 16445
rect 4433 16405 4445 16439
rect 4479 16405 4491 16439
rect 4433 16399 4491 16405
rect 4982 16396 4988 16448
rect 5040 16436 5046 16448
rect 5442 16436 5448 16448
rect 5040 16408 5448 16436
rect 5040 16396 5046 16408
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 5534 16396 5540 16448
rect 5592 16436 5598 16448
rect 5905 16439 5963 16445
rect 5905 16436 5917 16439
rect 5592 16408 5917 16436
rect 5592 16396 5598 16408
rect 5905 16405 5917 16408
rect 5951 16405 5963 16439
rect 5905 16399 5963 16405
rect 6086 16396 6092 16448
rect 6144 16436 6150 16448
rect 6748 16436 6776 16476
rect 6144 16408 6776 16436
rect 6144 16396 6150 16408
rect 6822 16396 6828 16448
rect 6880 16396 6886 16448
rect 8588 16445 8616 16476
rect 9030 16464 9036 16516
rect 9088 16504 9094 16516
rect 9398 16504 9404 16516
rect 9088 16476 9404 16504
rect 9088 16464 9094 16476
rect 9398 16464 9404 16476
rect 9456 16504 9462 16516
rect 11072 16504 11100 16535
rect 11238 16532 11244 16544
rect 11296 16532 11302 16584
rect 12894 16532 12900 16584
rect 12952 16532 12958 16584
rect 13078 16532 13084 16584
rect 13136 16532 13142 16584
rect 13170 16532 13176 16584
rect 13228 16572 13234 16584
rect 13265 16575 13323 16581
rect 13265 16572 13277 16575
rect 13228 16544 13277 16572
rect 13228 16532 13234 16544
rect 13265 16541 13277 16544
rect 13311 16572 13323 16575
rect 13556 16572 13584 16612
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 14921 16643 14979 16649
rect 14921 16609 14933 16643
rect 14967 16640 14979 16643
rect 15838 16640 15844 16652
rect 14967 16612 15844 16640
rect 14967 16609 14979 16612
rect 14921 16603 14979 16609
rect 15838 16600 15844 16612
rect 15896 16600 15902 16652
rect 13311 16544 13584 16572
rect 13311 16541 13323 16544
rect 13265 16535 13323 16541
rect 13630 16532 13636 16584
rect 13688 16532 13694 16584
rect 13722 16532 13728 16584
rect 13780 16572 13786 16584
rect 13817 16575 13875 16581
rect 13817 16572 13829 16575
rect 13780 16544 13829 16572
rect 13780 16532 13786 16544
rect 13817 16541 13829 16544
rect 13863 16541 13875 16575
rect 13817 16535 13875 16541
rect 15013 16575 15071 16581
rect 15013 16541 15025 16575
rect 15059 16541 15071 16575
rect 15013 16535 15071 16541
rect 15749 16575 15807 16581
rect 15749 16541 15761 16575
rect 15795 16572 15807 16575
rect 16022 16572 16028 16584
rect 15795 16544 16028 16572
rect 15795 16541 15807 16544
rect 15749 16535 15807 16541
rect 9456 16476 11100 16504
rect 9456 16464 9462 16476
rect 12434 16464 12440 16516
rect 12492 16504 12498 16516
rect 14826 16504 14832 16516
rect 12492 16476 14832 16504
rect 12492 16464 12498 16476
rect 14826 16464 14832 16476
rect 14884 16504 14890 16516
rect 15028 16504 15056 16535
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 16206 16532 16212 16584
rect 16264 16532 16270 16584
rect 16482 16532 16488 16584
rect 16540 16532 16546 16584
rect 16574 16532 16580 16584
rect 16632 16532 16638 16584
rect 15841 16507 15899 16513
rect 15841 16504 15853 16507
rect 14884 16476 15853 16504
rect 14884 16464 14890 16476
rect 15841 16473 15853 16476
rect 15887 16473 15899 16507
rect 15841 16467 15899 16473
rect 8573 16439 8631 16445
rect 8573 16405 8585 16439
rect 8619 16405 8631 16439
rect 8573 16399 8631 16405
rect 9122 16396 9128 16448
rect 9180 16396 9186 16448
rect 10226 16396 10232 16448
rect 10284 16436 10290 16448
rect 10597 16439 10655 16445
rect 10597 16436 10609 16439
rect 10284 16408 10609 16436
rect 10284 16396 10290 16408
rect 10597 16405 10609 16408
rect 10643 16405 10655 16439
rect 10597 16399 10655 16405
rect 13446 16396 13452 16448
rect 13504 16436 13510 16448
rect 13722 16436 13728 16448
rect 13504 16408 13728 16436
rect 13504 16396 13510 16408
rect 13722 16396 13728 16408
rect 13780 16396 13786 16448
rect 13906 16396 13912 16448
rect 13964 16436 13970 16448
rect 14691 16439 14749 16445
rect 14691 16436 14703 16439
rect 13964 16408 14703 16436
rect 13964 16396 13970 16408
rect 14691 16405 14703 16408
rect 14737 16436 14749 16439
rect 16758 16436 16764 16448
rect 14737 16408 16764 16436
rect 14737 16405 14749 16408
rect 14691 16399 14749 16405
rect 16758 16396 16764 16408
rect 16816 16396 16822 16448
rect 1104 16346 18400 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 18400 16346
rect 1104 16272 18400 16294
rect 5258 16232 5264 16244
rect 4816 16204 5264 16232
rect 2792 16136 4292 16164
rect 2590 16056 2596 16108
rect 2648 16096 2654 16108
rect 2792 16105 2820 16136
rect 2777 16099 2835 16105
rect 2777 16096 2789 16099
rect 2648 16068 2789 16096
rect 2648 16056 2654 16068
rect 2777 16065 2789 16068
rect 2823 16065 2835 16099
rect 2777 16059 2835 16065
rect 3050 16056 3056 16108
rect 3108 16096 3114 16108
rect 3145 16099 3203 16105
rect 3145 16096 3157 16099
rect 3108 16068 3157 16096
rect 3108 16056 3114 16068
rect 3145 16065 3157 16068
rect 3191 16065 3203 16099
rect 3145 16059 3203 16065
rect 4264 16028 4292 16136
rect 4816 16108 4844 16204
rect 5258 16192 5264 16204
rect 5316 16232 5322 16244
rect 5316 16204 5580 16232
rect 5316 16192 5322 16204
rect 5350 16124 5356 16176
rect 5408 16164 5414 16176
rect 5552 16164 5580 16204
rect 5626 16192 5632 16244
rect 5684 16192 5690 16244
rect 6917 16235 6975 16241
rect 6917 16232 6929 16235
rect 5752 16204 6929 16232
rect 5752 16164 5780 16204
rect 6917 16201 6929 16204
rect 6963 16232 6975 16235
rect 7653 16235 7711 16241
rect 7653 16232 7665 16235
rect 6963 16204 7665 16232
rect 6963 16201 6975 16204
rect 6917 16195 6975 16201
rect 7653 16201 7665 16204
rect 7699 16232 7711 16235
rect 7834 16232 7840 16244
rect 7699 16204 7840 16232
rect 7699 16201 7711 16204
rect 7653 16195 7711 16201
rect 7834 16192 7840 16204
rect 7892 16192 7898 16244
rect 7926 16192 7932 16244
rect 7984 16232 7990 16244
rect 8297 16235 8355 16241
rect 8297 16232 8309 16235
rect 7984 16204 8309 16232
rect 7984 16192 7990 16204
rect 8297 16201 8309 16204
rect 8343 16232 8355 16235
rect 8665 16235 8723 16241
rect 8665 16232 8677 16235
rect 8343 16204 8677 16232
rect 8343 16201 8355 16204
rect 8297 16195 8355 16201
rect 8665 16201 8677 16204
rect 8711 16201 8723 16235
rect 8665 16195 8723 16201
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 11149 16235 11207 16241
rect 11149 16232 11161 16235
rect 11112 16204 11161 16232
rect 11112 16192 11118 16204
rect 11149 16201 11161 16204
rect 11195 16232 11207 16235
rect 14274 16232 14280 16244
rect 11195 16204 14280 16232
rect 11195 16201 11207 16204
rect 11149 16195 11207 16201
rect 14274 16192 14280 16204
rect 14332 16192 14338 16244
rect 15838 16192 15844 16244
rect 15896 16192 15902 16244
rect 5408 16136 5488 16164
rect 5552 16136 5780 16164
rect 5408 16124 5414 16136
rect 4798 16056 4804 16108
rect 4856 16056 4862 16108
rect 5460 16096 5488 16136
rect 5644 16105 5672 16136
rect 5810 16124 5816 16176
rect 5868 16164 5874 16176
rect 6517 16167 6575 16173
rect 6517 16164 6529 16167
rect 5868 16136 6529 16164
rect 5868 16124 5874 16136
rect 6517 16133 6529 16136
rect 6563 16133 6575 16167
rect 6517 16127 6575 16133
rect 6730 16124 6736 16176
rect 6788 16164 6794 16176
rect 8113 16167 8171 16173
rect 8113 16164 8125 16167
rect 6788 16136 8125 16164
rect 6788 16124 6794 16136
rect 8113 16133 8125 16136
rect 8159 16133 8171 16167
rect 9030 16164 9036 16176
rect 8113 16127 8171 16133
rect 8588 16136 9036 16164
rect 5629 16099 5687 16105
rect 4908 16068 5396 16096
rect 5460 16068 5580 16096
rect 4908 16028 4936 16068
rect 4264 16000 4936 16028
rect 5074 15988 5080 16040
rect 5132 15988 5138 16040
rect 5166 15988 5172 16040
rect 5224 15988 5230 16040
rect 5258 15988 5264 16040
rect 5316 15988 5322 16040
rect 5368 16037 5396 16068
rect 5552 16037 5580 16068
rect 5629 16065 5641 16099
rect 5675 16065 5687 16099
rect 5629 16059 5687 16065
rect 5994 16056 6000 16108
rect 6052 16096 6058 16108
rect 6089 16099 6147 16105
rect 6089 16096 6101 16099
rect 6052 16068 6101 16096
rect 6052 16056 6058 16068
rect 6089 16065 6101 16068
rect 6135 16065 6147 16099
rect 6089 16059 6147 16065
rect 6822 16056 6828 16108
rect 6880 16056 6886 16108
rect 7101 16099 7159 16105
rect 7101 16065 7113 16099
rect 7147 16065 7159 16099
rect 7101 16059 7159 16065
rect 7193 16099 7251 16105
rect 7193 16065 7205 16099
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 7377 16099 7435 16105
rect 7377 16065 7389 16099
rect 7423 16065 7435 16099
rect 7377 16059 7435 16065
rect 7469 16099 7527 16105
rect 7469 16065 7481 16099
rect 7515 16065 7527 16099
rect 7469 16059 7527 16065
rect 5353 16031 5411 16037
rect 5353 15997 5365 16031
rect 5399 15997 5411 16031
rect 5353 15991 5411 15997
rect 5537 16031 5595 16037
rect 5537 15997 5549 16031
rect 5583 15997 5595 16031
rect 5813 16031 5871 16037
rect 5813 16028 5825 16031
rect 5537 15991 5595 15997
rect 5644 16000 5825 16028
rect 3326 15920 3332 15972
rect 3384 15960 3390 15972
rect 5092 15960 5120 15988
rect 3384 15932 5120 15960
rect 3384 15920 3390 15932
rect 4433 15895 4491 15901
rect 4433 15861 4445 15895
rect 4479 15892 4491 15895
rect 5258 15892 5264 15904
rect 4479 15864 5264 15892
rect 4479 15861 4491 15864
rect 4433 15855 4491 15861
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 5368 15892 5396 15991
rect 5442 15920 5448 15972
rect 5500 15960 5506 15972
rect 5644 15960 5672 16000
rect 5813 15997 5825 16000
rect 5859 16028 5871 16031
rect 7116 16028 7144 16059
rect 5859 16000 7144 16028
rect 5859 15997 5871 16000
rect 5813 15991 5871 15997
rect 5500 15932 5672 15960
rect 5500 15920 5506 15932
rect 5718 15920 5724 15972
rect 5776 15960 5782 15972
rect 5951 15963 6009 15969
rect 5951 15960 5963 15963
rect 5776 15932 5963 15960
rect 5776 15920 5782 15932
rect 5951 15929 5963 15932
rect 5997 15929 6009 15963
rect 5951 15923 6009 15929
rect 6380 15932 7052 15960
rect 5810 15892 5816 15904
rect 5368 15864 5816 15892
rect 5810 15852 5816 15864
rect 5868 15852 5874 15904
rect 6270 15852 6276 15904
rect 6328 15892 6334 15904
rect 6380 15901 6408 15932
rect 6365 15895 6423 15901
rect 6365 15892 6377 15895
rect 6328 15864 6377 15892
rect 6328 15852 6334 15864
rect 6365 15861 6377 15864
rect 6411 15861 6423 15895
rect 6365 15855 6423 15861
rect 6546 15852 6552 15904
rect 6604 15852 6610 15904
rect 7024 15892 7052 15932
rect 7098 15920 7104 15972
rect 7156 15920 7162 15972
rect 7208 15892 7236 16059
rect 7282 15988 7288 16040
rect 7340 15988 7346 16040
rect 7392 15960 7420 16059
rect 7484 16028 7512 16059
rect 7834 16056 7840 16108
rect 7892 16096 7898 16108
rect 7929 16099 7987 16105
rect 7929 16096 7941 16099
rect 7892 16068 7941 16096
rect 7892 16056 7898 16068
rect 7929 16065 7941 16068
rect 7975 16065 7987 16099
rect 8128 16096 8156 16127
rect 8294 16096 8300 16108
rect 8128 16068 8300 16096
rect 7929 16059 7987 16065
rect 8294 16056 8300 16068
rect 8352 16056 8358 16108
rect 8588 16105 8616 16136
rect 9030 16124 9036 16136
rect 9088 16164 9094 16176
rect 9861 16167 9919 16173
rect 9861 16164 9873 16167
rect 9088 16136 9873 16164
rect 9088 16124 9094 16136
rect 9861 16133 9873 16136
rect 9907 16133 9919 16167
rect 11885 16167 11943 16173
rect 11885 16164 11897 16167
rect 9861 16127 9919 16133
rect 11256 16136 11897 16164
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16065 8631 16099
rect 8573 16059 8631 16065
rect 8846 16056 8852 16108
rect 8904 16056 8910 16108
rect 9306 16056 9312 16108
rect 9364 16056 9370 16108
rect 9674 16056 9680 16108
rect 9732 16096 9738 16108
rect 10045 16099 10103 16105
rect 10045 16096 10057 16099
rect 9732 16068 10057 16096
rect 9732 16056 9738 16068
rect 10045 16065 10057 16068
rect 10091 16065 10103 16099
rect 10045 16059 10103 16065
rect 10134 16056 10140 16108
rect 10192 16096 10198 16108
rect 10689 16099 10747 16105
rect 10689 16096 10701 16099
rect 10192 16068 10701 16096
rect 10192 16056 10198 16068
rect 10689 16065 10701 16068
rect 10735 16065 10747 16099
rect 10689 16059 10747 16065
rect 11054 16056 11060 16108
rect 11112 16056 11118 16108
rect 11256 16105 11284 16136
rect 11241 16099 11299 16105
rect 11241 16065 11253 16099
rect 11287 16065 11299 16099
rect 11241 16059 11299 16065
rect 11330 16056 11336 16108
rect 11388 16096 11394 16108
rect 11716 16105 11744 16136
rect 11885 16133 11897 16136
rect 11931 16133 11943 16167
rect 11885 16127 11943 16133
rect 12066 16124 12072 16176
rect 12124 16124 12130 16176
rect 12250 16124 12256 16176
rect 12308 16124 12314 16176
rect 12434 16124 12440 16176
rect 12492 16124 12498 16176
rect 12526 16124 12532 16176
rect 12584 16164 12590 16176
rect 12897 16167 12955 16173
rect 12897 16164 12909 16167
rect 12584 16136 12909 16164
rect 12584 16124 12590 16136
rect 12897 16133 12909 16136
rect 12943 16133 12955 16167
rect 12897 16127 12955 16133
rect 13078 16124 13084 16176
rect 13136 16164 13142 16176
rect 13541 16167 13599 16173
rect 13541 16164 13553 16167
rect 13136 16136 13553 16164
rect 13136 16124 13142 16136
rect 13541 16133 13553 16136
rect 13587 16164 13599 16167
rect 13630 16164 13636 16176
rect 13587 16136 13636 16164
rect 13587 16133 13599 16136
rect 13541 16127 13599 16133
rect 13630 16124 13636 16136
rect 13688 16124 13694 16176
rect 16025 16167 16083 16173
rect 16025 16164 16037 16167
rect 15594 16136 16037 16164
rect 16025 16133 16037 16136
rect 16071 16133 16083 16167
rect 16025 16127 16083 16133
rect 16482 16124 16488 16176
rect 16540 16164 16546 16176
rect 17129 16167 17187 16173
rect 17129 16164 17141 16167
rect 16540 16136 17141 16164
rect 16540 16124 16546 16136
rect 17129 16133 17141 16136
rect 17175 16133 17187 16167
rect 17129 16127 17187 16133
rect 11517 16099 11575 16105
rect 11517 16096 11529 16099
rect 11388 16068 11529 16096
rect 11388 16056 11394 16068
rect 11517 16065 11529 16068
rect 11563 16065 11575 16099
rect 11517 16059 11575 16065
rect 11701 16099 11759 16105
rect 11701 16065 11713 16099
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 11793 16099 11851 16105
rect 11793 16065 11805 16099
rect 11839 16065 11851 16099
rect 11793 16059 11851 16065
rect 11977 16099 12035 16105
rect 11977 16065 11989 16099
rect 12023 16096 12035 16099
rect 12158 16096 12164 16108
rect 12023 16068 12164 16096
rect 12023 16065 12035 16068
rect 11977 16059 12035 16065
rect 8662 16028 8668 16040
rect 7484 16000 8668 16028
rect 8662 15988 8668 16000
rect 8720 16028 8726 16040
rect 8864 16028 8892 16056
rect 8720 16000 8892 16028
rect 8720 15988 8726 16000
rect 9582 15988 9588 16040
rect 9640 15988 9646 16040
rect 10229 16031 10287 16037
rect 10229 16028 10241 16031
rect 10152 16000 10241 16028
rect 7558 15960 7564 15972
rect 7392 15932 7564 15960
rect 7558 15920 7564 15932
rect 7616 15920 7622 15972
rect 7834 15920 7840 15972
rect 7892 15960 7898 15972
rect 9490 15960 9496 15972
rect 7892 15932 9496 15960
rect 7892 15920 7898 15932
rect 9490 15920 9496 15932
rect 9548 15920 9554 15972
rect 7024 15864 7236 15892
rect 8938 15852 8944 15904
rect 8996 15892 9002 15904
rect 9033 15895 9091 15901
rect 9033 15892 9045 15895
rect 8996 15864 9045 15892
rect 8996 15852 9002 15864
rect 9033 15861 9045 15864
rect 9079 15861 9091 15895
rect 9033 15855 9091 15861
rect 9122 15852 9128 15904
rect 9180 15892 9186 15904
rect 10152 15892 10180 16000
rect 10229 15997 10241 16000
rect 10275 16028 10287 16031
rect 10502 16028 10508 16040
rect 10275 16000 10508 16028
rect 10275 15997 10287 16000
rect 10229 15991 10287 15997
rect 10502 15988 10508 16000
rect 10560 15988 10566 16040
rect 10965 16031 11023 16037
rect 10965 15997 10977 16031
rect 11011 15997 11023 16031
rect 11808 16028 11836 16059
rect 12158 16056 12164 16068
rect 12216 16096 12222 16108
rect 12713 16099 12771 16105
rect 12713 16096 12725 16099
rect 12216 16068 12725 16096
rect 12216 16056 12222 16068
rect 12713 16065 12725 16068
rect 12759 16065 12771 16099
rect 12713 16059 12771 16065
rect 12805 16099 12863 16105
rect 12805 16065 12817 16099
rect 12851 16065 12863 16099
rect 12805 16059 12863 16065
rect 13357 16099 13415 16105
rect 13357 16065 13369 16099
rect 13403 16096 13415 16099
rect 13722 16096 13728 16108
rect 13403 16068 13728 16096
rect 13403 16065 13415 16068
rect 13357 16059 13415 16065
rect 12820 16028 12848 16059
rect 13722 16056 13728 16068
rect 13780 16056 13786 16108
rect 13814 16056 13820 16108
rect 13872 16056 13878 16108
rect 14090 16056 14096 16108
rect 14148 16056 14154 16108
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 16574 16096 16580 16108
rect 16163 16068 16580 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 16574 16056 16580 16068
rect 16632 16096 16638 16108
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 16632 16068 16865 16096
rect 16632 16056 16638 16068
rect 16853 16065 16865 16068
rect 16899 16096 16911 16099
rect 17034 16096 17040 16108
rect 16899 16068 17040 16096
rect 16899 16065 16911 16068
rect 16853 16059 16911 16065
rect 17034 16056 17040 16068
rect 17092 16056 17098 16108
rect 13078 16028 13084 16040
rect 11808 16000 13084 16028
rect 10965 15991 11023 15997
rect 10778 15920 10784 15972
rect 10836 15920 10842 15972
rect 10980 15960 11008 15991
rect 13078 15988 13084 16000
rect 13136 15988 13142 16040
rect 13173 16031 13231 16037
rect 13173 15997 13185 16031
rect 13219 16028 13231 16031
rect 13630 16028 13636 16040
rect 13219 16000 13636 16028
rect 13219 15997 13231 16000
rect 13173 15991 13231 15997
rect 13630 15988 13636 16000
rect 13688 15988 13694 16040
rect 14001 16031 14059 16037
rect 14001 15997 14013 16031
rect 14047 16028 14059 16031
rect 14369 16031 14427 16037
rect 14369 16028 14381 16031
rect 14047 16000 14381 16028
rect 14047 15997 14059 16000
rect 14001 15991 14059 15997
rect 14369 15997 14381 16000
rect 14415 15997 14427 16031
rect 14369 15991 14427 15997
rect 12529 15963 12587 15969
rect 12529 15960 12541 15963
rect 10980 15932 12541 15960
rect 12529 15929 12541 15932
rect 12575 15960 12587 15963
rect 13446 15960 13452 15972
rect 12575 15932 13452 15960
rect 12575 15929 12587 15932
rect 12529 15923 12587 15929
rect 13446 15920 13452 15932
rect 13504 15920 13510 15972
rect 9180 15864 10180 15892
rect 10873 15895 10931 15901
rect 9180 15852 9186 15864
rect 10873 15861 10885 15895
rect 10919 15892 10931 15895
rect 11054 15892 11060 15904
rect 10919 15864 11060 15892
rect 10919 15861 10931 15864
rect 10873 15855 10931 15861
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 11606 15852 11612 15904
rect 11664 15852 11670 15904
rect 16666 15852 16672 15904
rect 16724 15892 16730 15904
rect 16761 15895 16819 15901
rect 16761 15892 16773 15895
rect 16724 15864 16773 15892
rect 16724 15852 16730 15864
rect 16761 15861 16773 15864
rect 16807 15861 16819 15895
rect 16761 15855 16819 15861
rect 17126 15852 17132 15904
rect 17184 15892 17190 15904
rect 17221 15895 17279 15901
rect 17221 15892 17233 15895
rect 17184 15864 17233 15892
rect 17184 15852 17190 15864
rect 17221 15861 17233 15864
rect 17267 15861 17279 15895
rect 17221 15855 17279 15861
rect 1104 15802 18400 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 18400 15802
rect 1104 15728 18400 15750
rect 2685 15691 2743 15697
rect 2685 15657 2697 15691
rect 2731 15688 2743 15691
rect 2958 15688 2964 15700
rect 2731 15660 2964 15688
rect 2731 15657 2743 15660
rect 2685 15651 2743 15657
rect 2958 15648 2964 15660
rect 3016 15648 3022 15700
rect 3050 15648 3056 15700
rect 3108 15688 3114 15700
rect 3237 15691 3295 15697
rect 3237 15688 3249 15691
rect 3108 15660 3249 15688
rect 3108 15648 3114 15660
rect 3237 15657 3249 15660
rect 3283 15657 3295 15691
rect 3237 15651 3295 15657
rect 4522 15648 4528 15700
rect 4580 15688 4586 15700
rect 5994 15688 6000 15700
rect 4580 15660 6000 15688
rect 4580 15648 4586 15660
rect 5994 15648 6000 15660
rect 6052 15648 6058 15700
rect 6546 15648 6552 15700
rect 6604 15688 6610 15700
rect 9674 15688 9680 15700
rect 6604 15660 9680 15688
rect 6604 15648 6610 15660
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 9858 15688 9864 15700
rect 9784 15660 9864 15688
rect 2869 15623 2927 15629
rect 2869 15589 2881 15623
rect 2915 15620 2927 15623
rect 3326 15620 3332 15632
rect 2915 15592 3332 15620
rect 2915 15589 2927 15592
rect 2869 15583 2927 15589
rect 3326 15580 3332 15592
rect 3384 15580 3390 15632
rect 6730 15620 6736 15632
rect 4908 15592 6736 15620
rect 3510 15552 3516 15564
rect 2516 15524 3516 15552
rect 2516 15493 2544 15524
rect 3510 15512 3516 15524
rect 3568 15512 3574 15564
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15552 4491 15555
rect 4614 15552 4620 15564
rect 4479 15524 4620 15552
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 4614 15512 4620 15524
rect 4672 15512 4678 15564
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15453 2559 15487
rect 2501 15447 2559 15453
rect 2590 15444 2596 15496
rect 2648 15484 2654 15496
rect 2685 15487 2743 15493
rect 2685 15484 2697 15487
rect 2648 15456 2697 15484
rect 2648 15444 2654 15456
rect 2685 15453 2697 15456
rect 2731 15484 2743 15487
rect 4249 15487 4307 15493
rect 2731 15456 3280 15484
rect 2731 15453 2743 15456
rect 2685 15447 2743 15453
rect 3252 15425 3280 15456
rect 4249 15453 4261 15487
rect 4295 15484 4307 15487
rect 4798 15484 4804 15496
rect 4295 15456 4804 15484
rect 4295 15453 4307 15456
rect 4249 15447 4307 15453
rect 4798 15444 4804 15456
rect 4856 15444 4862 15496
rect 4908 15493 4936 15592
rect 6730 15580 6736 15592
rect 6788 15580 6794 15632
rect 8018 15580 8024 15632
rect 8076 15620 8082 15632
rect 9125 15623 9183 15629
rect 9125 15620 9137 15623
rect 8076 15592 9137 15620
rect 8076 15580 8082 15592
rect 9125 15589 9137 15592
rect 9171 15620 9183 15623
rect 9784 15620 9812 15660
rect 9858 15648 9864 15660
rect 9916 15648 9922 15700
rect 9950 15648 9956 15700
rect 10008 15648 10014 15700
rect 11698 15648 11704 15700
rect 11756 15688 11762 15700
rect 15105 15691 15163 15697
rect 15105 15688 15117 15691
rect 11756 15660 15117 15688
rect 11756 15648 11762 15660
rect 15105 15657 15117 15660
rect 15151 15688 15163 15691
rect 15746 15688 15752 15700
rect 15151 15660 15752 15688
rect 15151 15657 15163 15660
rect 15105 15651 15163 15657
rect 15746 15648 15752 15660
rect 15804 15648 15810 15700
rect 17770 15620 17776 15632
rect 9171 15592 9812 15620
rect 17144 15592 17776 15620
rect 9171 15589 9183 15592
rect 9125 15583 9183 15589
rect 4985 15555 5043 15561
rect 4985 15521 4997 15555
rect 5031 15521 5043 15555
rect 6270 15552 6276 15564
rect 4985 15515 5043 15521
rect 5185 15524 6276 15552
rect 4893 15487 4951 15493
rect 4893 15453 4905 15487
rect 4939 15453 4951 15487
rect 4893 15447 4951 15453
rect 3237 15419 3295 15425
rect 3237 15385 3249 15419
rect 3283 15385 3295 15419
rect 4430 15416 4436 15428
rect 3237 15379 3295 15385
rect 3436 15388 4436 15416
rect 3436 15357 3464 15388
rect 4430 15376 4436 15388
rect 4488 15416 4494 15428
rect 4525 15419 4583 15425
rect 4525 15416 4537 15419
rect 4488 15388 4537 15416
rect 4488 15376 4494 15388
rect 4525 15385 4537 15388
rect 4571 15416 4583 15419
rect 4706 15416 4712 15428
rect 4571 15388 4712 15416
rect 4571 15385 4583 15388
rect 4525 15379 4583 15385
rect 4706 15376 4712 15388
rect 4764 15376 4770 15428
rect 5000 15416 5028 15515
rect 5185 15493 5213 15524
rect 6270 15512 6276 15524
rect 6328 15512 6334 15564
rect 8573 15555 8631 15561
rect 8573 15552 8585 15555
rect 8128 15524 8585 15552
rect 5169 15487 5227 15493
rect 5169 15453 5181 15487
rect 5215 15453 5227 15487
rect 5169 15447 5227 15453
rect 5261 15487 5319 15493
rect 5261 15453 5273 15487
rect 5307 15453 5319 15487
rect 5534 15484 5540 15496
rect 5261 15447 5319 15453
rect 5368 15456 5540 15484
rect 4908 15388 5028 15416
rect 3421 15351 3479 15357
rect 3421 15317 3433 15351
rect 3467 15317 3479 15351
rect 3421 15311 3479 15317
rect 4065 15351 4123 15357
rect 4065 15317 4077 15351
rect 4111 15348 4123 15351
rect 4246 15348 4252 15360
rect 4111 15320 4252 15348
rect 4111 15317 4123 15320
rect 4065 15311 4123 15317
rect 4246 15308 4252 15320
rect 4304 15308 4310 15360
rect 4614 15308 4620 15360
rect 4672 15348 4678 15360
rect 4908 15348 4936 15388
rect 5074 15376 5080 15428
rect 5132 15416 5138 15428
rect 5276 15416 5304 15447
rect 5132 15388 5304 15416
rect 5132 15376 5138 15388
rect 4672 15320 4936 15348
rect 4672 15308 4678 15320
rect 5166 15308 5172 15360
rect 5224 15348 5230 15360
rect 5368 15348 5396 15456
rect 5534 15444 5540 15456
rect 5592 15444 5598 15496
rect 5810 15444 5816 15496
rect 5868 15484 5874 15496
rect 5905 15487 5963 15493
rect 5905 15484 5917 15487
rect 5868 15456 5917 15484
rect 5868 15444 5874 15456
rect 5905 15453 5917 15456
rect 5951 15453 5963 15487
rect 5905 15447 5963 15453
rect 6457 15487 6515 15493
rect 6457 15453 6469 15487
rect 6503 15484 6515 15487
rect 7558 15484 7564 15496
rect 6503 15456 7564 15484
rect 6503 15453 6515 15456
rect 6457 15447 6515 15453
rect 7558 15444 7564 15456
rect 7616 15444 7622 15496
rect 7742 15444 7748 15496
rect 7800 15444 7806 15496
rect 7926 15493 7932 15496
rect 7893 15487 7932 15493
rect 7893 15453 7905 15487
rect 7893 15447 7932 15453
rect 7926 15444 7932 15447
rect 7984 15444 7990 15496
rect 8128 15493 8156 15524
rect 8573 15521 8585 15524
rect 8619 15521 8631 15555
rect 8573 15515 8631 15521
rect 9030 15512 9036 15564
rect 9088 15512 9094 15564
rect 9674 15552 9680 15564
rect 9508 15524 9680 15552
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15453 8171 15487
rect 8113 15447 8171 15453
rect 8202 15444 8208 15496
rect 8260 15493 8266 15496
rect 8260 15484 8268 15493
rect 8665 15487 8723 15493
rect 8260 15456 8305 15484
rect 8260 15447 8268 15456
rect 8665 15453 8677 15487
rect 8711 15484 8723 15487
rect 8754 15484 8760 15496
rect 8711 15456 8760 15484
rect 8711 15453 8723 15456
rect 8665 15447 8723 15453
rect 8260 15444 8266 15447
rect 5445 15419 5503 15425
rect 5445 15385 5457 15419
rect 5491 15416 5503 15419
rect 5491 15388 5580 15416
rect 5491 15385 5503 15388
rect 5445 15379 5503 15385
rect 5224 15320 5396 15348
rect 5552 15348 5580 15388
rect 6086 15376 6092 15428
rect 6144 15416 6150 15428
rect 6641 15419 6699 15425
rect 6641 15416 6653 15419
rect 6144 15388 6653 15416
rect 6144 15376 6150 15388
rect 6641 15385 6653 15388
rect 6687 15385 6699 15419
rect 6641 15379 6699 15385
rect 6454 15348 6460 15360
rect 5552 15320 6460 15348
rect 5224 15308 5230 15320
rect 6454 15308 6460 15320
rect 6512 15308 6518 15360
rect 6656 15348 6684 15379
rect 7282 15376 7288 15428
rect 7340 15416 7346 15428
rect 8018 15416 8024 15428
rect 7340 15388 8024 15416
rect 7340 15376 7346 15388
rect 8018 15376 8024 15388
rect 8076 15376 8082 15428
rect 8680 15416 8708 15447
rect 8754 15444 8760 15456
rect 8812 15444 8818 15496
rect 9398 15444 9404 15496
rect 9456 15444 9462 15496
rect 9508 15493 9536 15524
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 15289 15555 15347 15561
rect 15289 15521 15301 15555
rect 15335 15552 15347 15555
rect 17144 15552 17172 15592
rect 17770 15580 17776 15592
rect 17828 15580 17834 15632
rect 15335 15524 17172 15552
rect 15335 15521 15347 15524
rect 15289 15515 15347 15521
rect 17218 15512 17224 15564
rect 17276 15512 17282 15564
rect 9493 15487 9551 15493
rect 9493 15453 9505 15487
rect 9539 15453 9551 15487
rect 9493 15447 9551 15453
rect 9582 15444 9588 15496
rect 9640 15484 9646 15496
rect 9766 15484 9772 15496
rect 9640 15456 9772 15484
rect 9640 15444 9646 15456
rect 9766 15444 9772 15456
rect 9824 15484 9830 15496
rect 9861 15487 9919 15493
rect 9861 15484 9873 15487
rect 9824 15456 9873 15484
rect 9824 15444 9830 15456
rect 9861 15453 9873 15456
rect 9907 15453 9919 15487
rect 9861 15447 9919 15453
rect 9953 15487 10011 15493
rect 9953 15453 9965 15487
rect 9999 15484 10011 15487
rect 9999 15456 10088 15484
rect 9999 15453 10011 15456
rect 9953 15447 10011 15453
rect 10060 15428 10088 15456
rect 12618 15444 12624 15496
rect 12676 15484 12682 15496
rect 12713 15487 12771 15493
rect 12713 15484 12725 15487
rect 12676 15456 12725 15484
rect 12676 15444 12682 15456
rect 12713 15453 12725 15456
rect 12759 15453 12771 15487
rect 12713 15447 12771 15453
rect 8128 15388 8708 15416
rect 8128 15348 8156 15388
rect 9306 15376 9312 15428
rect 9364 15376 9370 15428
rect 10042 15376 10048 15428
rect 10100 15376 10106 15428
rect 10686 15376 10692 15428
rect 10744 15416 10750 15428
rect 12434 15416 12440 15428
rect 10744 15388 12440 15416
rect 10744 15376 10750 15388
rect 12434 15376 12440 15388
rect 12492 15376 12498 15428
rect 12728 15416 12756 15447
rect 14918 15444 14924 15496
rect 14976 15444 14982 15496
rect 16666 15444 16672 15496
rect 16724 15444 16730 15496
rect 16850 15444 16856 15496
rect 16908 15484 16914 15496
rect 17129 15487 17187 15493
rect 17129 15484 17141 15487
rect 16908 15456 17141 15484
rect 16908 15444 16914 15456
rect 17129 15453 17141 15456
rect 17175 15453 17187 15487
rect 17129 15447 17187 15453
rect 17494 15444 17500 15496
rect 17552 15493 17558 15496
rect 17552 15487 17589 15493
rect 17577 15453 17589 15487
rect 17552 15447 17589 15453
rect 17552 15444 17558 15447
rect 12728 15388 14964 15416
rect 6656 15320 8156 15348
rect 8386 15308 8392 15360
rect 8444 15308 8450 15360
rect 9769 15351 9827 15357
rect 9769 15317 9781 15351
rect 9815 15348 9827 15351
rect 9858 15348 9864 15360
rect 9815 15320 9864 15348
rect 9815 15317 9827 15320
rect 9769 15311 9827 15317
rect 9858 15308 9864 15320
rect 9916 15308 9922 15360
rect 9950 15308 9956 15360
rect 10008 15348 10014 15360
rect 10229 15351 10287 15357
rect 10229 15348 10241 15351
rect 10008 15320 10241 15348
rect 10008 15308 10014 15320
rect 10229 15317 10241 15320
rect 10275 15317 10287 15351
rect 10229 15311 10287 15317
rect 10778 15308 10784 15360
rect 10836 15348 10842 15360
rect 12158 15348 12164 15360
rect 10836 15320 12164 15348
rect 10836 15308 10842 15320
rect 12158 15308 12164 15320
rect 12216 15348 12222 15360
rect 12897 15351 12955 15357
rect 12897 15348 12909 15351
rect 12216 15320 12909 15348
rect 12216 15308 12222 15320
rect 12897 15317 12909 15320
rect 12943 15348 12955 15351
rect 13170 15348 13176 15360
rect 12943 15320 13176 15348
rect 12943 15317 12955 15320
rect 12897 15311 12955 15317
rect 13170 15308 13176 15320
rect 13228 15308 13234 15360
rect 14936 15348 14964 15388
rect 15010 15376 15016 15428
rect 15068 15416 15074 15428
rect 15565 15419 15623 15425
rect 15565 15416 15577 15419
rect 15068 15388 15577 15416
rect 15068 15376 15074 15388
rect 15565 15385 15577 15388
rect 15611 15385 15623 15419
rect 15565 15379 15623 15385
rect 15930 15348 15936 15360
rect 14936 15320 15936 15348
rect 15930 15308 15936 15320
rect 15988 15308 15994 15360
rect 16574 15308 16580 15360
rect 16632 15348 16638 15360
rect 17037 15351 17095 15357
rect 17037 15348 17049 15351
rect 16632 15320 17049 15348
rect 16632 15308 16638 15320
rect 17037 15317 17049 15320
rect 17083 15317 17095 15351
rect 17037 15311 17095 15317
rect 17586 15308 17592 15360
rect 17644 15348 17650 15360
rect 17681 15351 17739 15357
rect 17681 15348 17693 15351
rect 17644 15320 17693 15348
rect 17644 15308 17650 15320
rect 17681 15317 17693 15320
rect 17727 15317 17739 15351
rect 17681 15311 17739 15317
rect 1104 15258 18400 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 18400 15258
rect 1104 15184 18400 15206
rect 4430 15104 4436 15156
rect 4488 15144 4494 15156
rect 5350 15144 5356 15156
rect 4488 15116 5356 15144
rect 4488 15104 4494 15116
rect 5350 15104 5356 15116
rect 5408 15104 5414 15156
rect 7374 15104 7380 15156
rect 7432 15144 7438 15156
rect 7745 15147 7803 15153
rect 7745 15144 7757 15147
rect 7432 15116 7757 15144
rect 7432 15104 7438 15116
rect 7745 15113 7757 15116
rect 7791 15113 7803 15147
rect 7745 15107 7803 15113
rect 7926 15104 7932 15156
rect 7984 15104 7990 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 8849 15147 8907 15153
rect 8849 15144 8861 15147
rect 8352 15116 8861 15144
rect 8352 15104 8358 15116
rect 8849 15113 8861 15116
rect 8895 15144 8907 15147
rect 10042 15144 10048 15156
rect 8895 15116 10048 15144
rect 8895 15113 8907 15116
rect 8849 15107 8907 15113
rect 10042 15104 10048 15116
rect 10100 15104 10106 15156
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 10796 15116 11529 15144
rect 3789 15079 3847 15085
rect 3789 15076 3801 15079
rect 2332 15048 3801 15076
rect 2038 14968 2044 15020
rect 2096 14968 2102 15020
rect 2332 15017 2360 15048
rect 3789 15045 3801 15048
rect 3835 15045 3847 15079
rect 5902 15076 5908 15088
rect 3789 15039 3847 15045
rect 5276 15048 5908 15076
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 14977 2375 15011
rect 2317 14971 2375 14977
rect 2406 14968 2412 15020
rect 2464 14968 2470 15020
rect 2498 14968 2504 15020
rect 2556 15008 2562 15020
rect 2593 15011 2651 15017
rect 2593 15008 2605 15011
rect 2556 14980 2605 15008
rect 2556 14968 2562 14980
rect 2593 14977 2605 14980
rect 2639 14977 2651 15011
rect 2593 14971 2651 14977
rect 2685 15011 2743 15017
rect 2685 14977 2697 15011
rect 2731 15008 2743 15011
rect 2866 15008 2872 15020
rect 2731 14980 2872 15008
rect 2731 14977 2743 14980
rect 2685 14971 2743 14977
rect 2866 14968 2872 14980
rect 2924 14968 2930 15020
rect 3053 15011 3111 15017
rect 3053 14977 3065 15011
rect 3099 15008 3111 15011
rect 3694 15008 3700 15020
rect 3099 14980 3700 15008
rect 3099 14977 3111 14980
rect 3053 14971 3111 14977
rect 3694 14968 3700 14980
rect 3752 14968 3758 15020
rect 3970 14968 3976 15020
rect 4028 14968 4034 15020
rect 4062 14968 4068 15020
rect 4120 15008 4126 15020
rect 4157 15011 4215 15017
rect 4157 15008 4169 15011
rect 4120 14980 4169 15008
rect 4120 14968 4126 14980
rect 4157 14977 4169 14980
rect 4203 14977 4215 15011
rect 4157 14971 4215 14977
rect 4246 14968 4252 15020
rect 4304 14968 4310 15020
rect 1765 14943 1823 14949
rect 1765 14909 1777 14943
rect 1811 14940 1823 14943
rect 2133 14943 2191 14949
rect 2133 14940 2145 14943
rect 1811 14912 2145 14940
rect 1811 14909 1823 14912
rect 1765 14903 1823 14909
rect 2133 14909 2145 14912
rect 2179 14909 2191 14943
rect 2424 14940 2452 14968
rect 2777 14943 2835 14949
rect 2777 14940 2789 14943
rect 2424 14912 2789 14940
rect 2133 14903 2191 14909
rect 2777 14909 2789 14912
rect 2823 14909 2835 14943
rect 2777 14903 2835 14909
rect 2958 14900 2964 14952
rect 3016 14900 3022 14952
rect 3145 14943 3203 14949
rect 3145 14909 3157 14943
rect 3191 14909 3203 14943
rect 3145 14903 3203 14909
rect 3160 14872 3188 14903
rect 3234 14900 3240 14952
rect 3292 14900 3298 14952
rect 5276 14872 5304 15048
rect 5902 15036 5908 15048
rect 5960 15036 5966 15088
rect 6822 15036 6828 15088
rect 6880 15076 6886 15088
rect 7285 15079 7343 15085
rect 7285 15076 7297 15079
rect 6880 15048 7297 15076
rect 6880 15036 6886 15048
rect 7285 15045 7297 15048
rect 7331 15045 7343 15079
rect 7944 15076 7972 15104
rect 7285 15039 7343 15045
rect 7392 15048 7972 15076
rect 7392 15020 7420 15048
rect 8018 15036 8024 15088
rect 8076 15076 8082 15088
rect 9398 15085 9404 15088
rect 9385 15079 9404 15085
rect 9385 15076 9397 15079
rect 8076 15048 9397 15076
rect 8076 15036 8082 15048
rect 9385 15045 9397 15048
rect 9385 15039 9404 15045
rect 9398 15036 9404 15039
rect 9456 15036 9462 15088
rect 9582 15036 9588 15088
rect 9640 15036 9646 15088
rect 9858 15036 9864 15088
rect 9916 15076 9922 15088
rect 9916 15048 10548 15076
rect 9916 15036 9922 15048
rect 5350 14968 5356 15020
rect 5408 15008 5414 15020
rect 5537 15011 5595 15017
rect 5537 15008 5549 15011
rect 5408 14980 5549 15008
rect 5408 14968 5414 14980
rect 5537 14977 5549 14980
rect 5583 14977 5595 15011
rect 5537 14971 5595 14977
rect 5721 15011 5779 15017
rect 5721 14977 5733 15011
rect 5767 14977 5779 15011
rect 5721 14971 5779 14977
rect 5736 14940 5764 14971
rect 7006 14968 7012 15020
rect 7064 15008 7070 15020
rect 7193 15011 7251 15017
rect 7193 15008 7205 15011
rect 7064 14980 7205 15008
rect 7064 14968 7070 14980
rect 7193 14977 7205 14980
rect 7239 14977 7251 15011
rect 7193 14971 7251 14977
rect 7374 14968 7380 15020
rect 7432 14968 7438 15020
rect 7558 14968 7564 15020
rect 7616 14968 7622 15020
rect 7653 15011 7711 15017
rect 7653 14977 7665 15011
rect 7699 15008 7711 15011
rect 7834 15008 7840 15020
rect 7699 14980 7840 15008
rect 7699 14977 7711 14980
rect 7653 14971 7711 14977
rect 7668 14940 7696 14971
rect 7834 14968 7840 14980
rect 7892 14968 7898 15020
rect 7926 14968 7932 15020
rect 7984 14968 7990 15020
rect 9033 15011 9091 15017
rect 9033 15008 9045 15011
rect 8036 14980 9045 15008
rect 5736 14912 7696 14940
rect 3160 14844 5304 14872
rect 5534 14832 5540 14884
rect 5592 14872 5598 14884
rect 8036 14872 8064 14980
rect 9033 14977 9045 14980
rect 9079 15008 9091 15011
rect 9953 15011 10011 15017
rect 9079 14980 9812 15008
rect 9079 14977 9091 14980
rect 9033 14971 9091 14977
rect 8113 14943 8171 14949
rect 8113 14909 8125 14943
rect 8159 14909 8171 14943
rect 8113 14903 8171 14909
rect 5592 14844 8064 14872
rect 5592 14832 5598 14844
rect 1670 14764 1676 14816
rect 1728 14804 1734 14816
rect 1857 14807 1915 14813
rect 1857 14804 1869 14807
rect 1728 14776 1869 14804
rect 1728 14764 1734 14776
rect 1857 14773 1869 14776
rect 1903 14773 1915 14807
rect 1857 14767 1915 14773
rect 1946 14764 1952 14816
rect 2004 14764 2010 14816
rect 2222 14764 2228 14816
rect 2280 14804 2286 14816
rect 3234 14804 3240 14816
rect 2280 14776 3240 14804
rect 2280 14764 2286 14776
rect 3234 14764 3240 14776
rect 3292 14764 3298 14816
rect 5905 14807 5963 14813
rect 5905 14773 5917 14807
rect 5951 14804 5963 14807
rect 6822 14804 6828 14816
rect 5951 14776 6828 14804
rect 5951 14773 5963 14776
rect 5905 14767 5963 14773
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7009 14807 7067 14813
rect 7009 14773 7021 14807
rect 7055 14804 7067 14807
rect 7282 14804 7288 14816
rect 7055 14776 7288 14804
rect 7055 14773 7067 14776
rect 7009 14767 7067 14773
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 7374 14764 7380 14816
rect 7432 14804 7438 14816
rect 7558 14804 7564 14816
rect 7432 14776 7564 14804
rect 7432 14764 7438 14776
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 7834 14764 7840 14816
rect 7892 14804 7898 14816
rect 8128 14804 8156 14903
rect 8202 14832 8208 14884
rect 8260 14872 8266 14884
rect 9784 14881 9812 14980
rect 9953 14977 9965 15011
rect 9999 14977 10011 15011
rect 9953 14971 10011 14977
rect 9968 14940 9996 14971
rect 10410 14968 10416 15020
rect 10468 14968 10474 15020
rect 10520 15017 10548 15048
rect 10686 15036 10692 15088
rect 10744 15036 10750 15088
rect 10796 15085 10824 15116
rect 11517 15113 11529 15116
rect 11563 15113 11575 15147
rect 11517 15107 11575 15113
rect 11974 15104 11980 15156
rect 12032 15144 12038 15156
rect 12345 15147 12403 15153
rect 12345 15144 12357 15147
rect 12032 15116 12357 15144
rect 12032 15104 12038 15116
rect 12345 15113 12357 15116
rect 12391 15113 12403 15147
rect 12345 15107 12403 15113
rect 15194 15104 15200 15156
rect 15252 15104 15258 15156
rect 15470 15104 15476 15156
rect 15528 15144 15534 15156
rect 16853 15147 16911 15153
rect 16853 15144 16865 15147
rect 15528 15116 16865 15144
rect 15528 15104 15534 15116
rect 16853 15113 16865 15116
rect 16899 15113 16911 15147
rect 16853 15107 16911 15113
rect 17034 15104 17040 15156
rect 17092 15144 17098 15156
rect 17218 15144 17224 15156
rect 17092 15116 17224 15144
rect 17092 15104 17098 15116
rect 17218 15104 17224 15116
rect 17276 15144 17282 15156
rect 17681 15147 17739 15153
rect 17681 15144 17693 15147
rect 17276 15116 17693 15144
rect 17276 15104 17282 15116
rect 17681 15113 17693 15116
rect 17727 15113 17739 15147
rect 17681 15107 17739 15113
rect 10781 15079 10839 15085
rect 10781 15045 10793 15079
rect 10827 15045 10839 15079
rect 10781 15039 10839 15045
rect 10962 15036 10968 15088
rect 11020 15076 11026 15088
rect 12250 15076 12256 15088
rect 11020 15048 12256 15076
rect 11020 15036 11026 15048
rect 12250 15036 12256 15048
rect 12308 15076 12314 15088
rect 12713 15079 12771 15085
rect 12713 15076 12725 15079
rect 12308 15048 12725 15076
rect 12308 15036 12314 15048
rect 12713 15045 12725 15048
rect 12759 15045 12771 15079
rect 12713 15039 12771 15045
rect 12802 15036 12808 15088
rect 12860 15085 12866 15088
rect 12860 15079 12889 15085
rect 12877 15045 12889 15079
rect 12860 15039 12889 15045
rect 16485 15079 16543 15085
rect 16485 15045 16497 15079
rect 16531 15076 16543 15079
rect 18046 15076 18052 15088
rect 16531 15048 18052 15076
rect 16531 15045 16543 15048
rect 16485 15039 16543 15045
rect 12860 15036 12866 15039
rect 18046 15036 18052 15048
rect 18104 15036 18110 15088
rect 10505 15011 10563 15017
rect 10505 14977 10517 15011
rect 10551 14977 10563 15011
rect 10505 14971 10563 14977
rect 10870 14968 10876 15020
rect 10928 14968 10934 15020
rect 11606 14968 11612 15020
rect 11664 15008 11670 15020
rect 12069 15011 12127 15017
rect 12069 15008 12081 15011
rect 11664 14980 12081 15008
rect 11664 14968 11670 14980
rect 12069 14977 12081 14980
rect 12115 14977 12127 15011
rect 12069 14971 12127 14977
rect 12526 14968 12532 15020
rect 12584 14968 12590 15020
rect 12621 15011 12679 15017
rect 12621 14977 12633 15011
rect 12667 15008 12679 15011
rect 12667 14980 12940 15008
rect 12667 14977 12679 14980
rect 12621 14971 12679 14977
rect 12912 14952 12940 14980
rect 13170 14968 13176 15020
rect 13228 15008 13234 15020
rect 13357 15011 13415 15017
rect 13357 15008 13369 15011
rect 13228 14980 13369 15008
rect 13228 14968 13234 14980
rect 13357 14977 13369 14980
rect 13403 14977 13415 15011
rect 13357 14971 13415 14977
rect 13446 14968 13452 15020
rect 13504 14968 13510 15020
rect 15746 14968 15752 15020
rect 15804 15008 15810 15020
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 15804 14980 16681 15008
rect 15804 14968 15810 14980
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 16942 14968 16948 15020
rect 17000 14968 17006 15020
rect 17037 15011 17095 15017
rect 17037 14977 17049 15011
rect 17083 15008 17095 15011
rect 17126 15008 17132 15020
rect 17083 14980 17132 15008
rect 17083 14977 17095 14980
rect 17037 14971 17095 14977
rect 17126 14968 17132 14980
rect 17184 14968 17190 15020
rect 17954 14968 17960 15020
rect 18012 14968 18018 15020
rect 11422 14940 11428 14952
rect 9968 14912 11428 14940
rect 11422 14900 11428 14912
rect 11480 14900 11486 14952
rect 11793 14943 11851 14949
rect 11793 14909 11805 14943
rect 11839 14940 11851 14943
rect 12802 14940 12808 14952
rect 11839 14912 12808 14940
rect 11839 14909 11851 14912
rect 11793 14903 11851 14909
rect 12802 14900 12808 14912
rect 12860 14900 12866 14952
rect 12894 14900 12900 14952
rect 12952 14900 12958 14952
rect 12986 14900 12992 14952
rect 13044 14900 13050 14952
rect 13078 14900 13084 14952
rect 13136 14940 13142 14952
rect 13265 14943 13323 14949
rect 13265 14940 13277 14943
rect 13136 14912 13277 14940
rect 13136 14900 13142 14912
rect 13265 14909 13277 14912
rect 13311 14909 13323 14943
rect 13265 14903 13323 14909
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14940 13599 14943
rect 13722 14940 13728 14952
rect 13587 14912 13728 14940
rect 13587 14909 13599 14912
rect 13541 14903 13599 14909
rect 9769 14875 9827 14881
rect 8260 14844 9536 14872
rect 8260 14832 8266 14844
rect 7892 14776 8156 14804
rect 7892 14764 7898 14776
rect 8938 14764 8944 14816
rect 8996 14804 9002 14816
rect 9217 14807 9275 14813
rect 9217 14804 9229 14807
rect 8996 14776 9229 14804
rect 8996 14764 9002 14776
rect 9217 14773 9229 14776
rect 9263 14773 9275 14807
rect 9217 14767 9275 14773
rect 9306 14764 9312 14816
rect 9364 14804 9370 14816
rect 9401 14807 9459 14813
rect 9401 14804 9413 14807
rect 9364 14776 9413 14804
rect 9364 14764 9370 14776
rect 9401 14773 9413 14776
rect 9447 14773 9459 14807
rect 9508 14804 9536 14844
rect 9769 14841 9781 14875
rect 9815 14841 9827 14875
rect 9769 14835 9827 14841
rect 11057 14875 11115 14881
rect 11057 14841 11069 14875
rect 11103 14872 11115 14875
rect 13280 14872 13308 14903
rect 13722 14900 13728 14912
rect 13780 14940 13786 14952
rect 14550 14940 14556 14952
rect 13780 14912 14556 14940
rect 13780 14900 13786 14912
rect 14550 14900 14556 14912
rect 14608 14900 14614 14952
rect 16298 14872 16304 14884
rect 11103 14844 13216 14872
rect 13280 14844 16304 14872
rect 11103 14841 11115 14844
rect 11057 14835 11115 14841
rect 11701 14807 11759 14813
rect 11701 14804 11713 14807
rect 9508 14776 11713 14804
rect 9401 14767 9459 14773
rect 11701 14773 11713 14776
rect 11747 14773 11759 14807
rect 11701 14767 11759 14773
rect 12710 14764 12716 14816
rect 12768 14804 12774 14816
rect 13081 14807 13139 14813
rect 13081 14804 13093 14807
rect 12768 14776 13093 14804
rect 12768 14764 12774 14776
rect 13081 14773 13093 14776
rect 13127 14773 13139 14807
rect 13188 14804 13216 14844
rect 16298 14832 16304 14844
rect 16356 14872 16362 14884
rect 17221 14875 17279 14881
rect 17221 14872 17233 14875
rect 16356 14844 17233 14872
rect 16356 14832 16362 14844
rect 17221 14841 17233 14844
rect 17267 14872 17279 14875
rect 17494 14872 17500 14884
rect 17267 14844 17500 14872
rect 17267 14841 17279 14844
rect 17221 14835 17279 14841
rect 17494 14832 17500 14844
rect 17552 14832 17558 14884
rect 15470 14804 15476 14816
rect 13188 14776 15476 14804
rect 13081 14767 13139 14773
rect 15470 14764 15476 14776
rect 15528 14764 15534 14816
rect 15654 14764 15660 14816
rect 15712 14804 15718 14816
rect 16669 14807 16727 14813
rect 16669 14804 16681 14807
rect 15712 14776 16681 14804
rect 15712 14764 15718 14776
rect 16669 14773 16681 14776
rect 16715 14773 16727 14807
rect 16669 14767 16727 14773
rect 1104 14714 18400 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 18400 14714
rect 1104 14640 18400 14662
rect 1946 14560 1952 14612
rect 2004 14600 2010 14612
rect 2317 14603 2375 14609
rect 2317 14600 2329 14603
rect 2004 14572 2329 14600
rect 2004 14560 2010 14572
rect 2317 14569 2329 14572
rect 2363 14569 2375 14603
rect 2317 14563 2375 14569
rect 2682 14560 2688 14612
rect 2740 14600 2746 14612
rect 6365 14603 6423 14609
rect 6365 14600 6377 14603
rect 2740 14572 6377 14600
rect 2740 14560 2746 14572
rect 6365 14569 6377 14572
rect 6411 14569 6423 14603
rect 6365 14563 6423 14569
rect 6454 14560 6460 14612
rect 6512 14560 6518 14612
rect 7193 14603 7251 14609
rect 7193 14569 7205 14603
rect 7239 14600 7251 14603
rect 7926 14600 7932 14612
rect 7239 14572 7932 14600
rect 7239 14569 7251 14572
rect 7193 14563 7251 14569
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 9122 14600 9128 14612
rect 8036 14572 9128 14600
rect 842 14492 848 14544
rect 900 14532 906 14544
rect 1489 14535 1547 14541
rect 1489 14532 1501 14535
rect 900 14504 1501 14532
rect 900 14492 906 14504
rect 1489 14501 1501 14504
rect 1535 14501 1547 14535
rect 1489 14495 1547 14501
rect 3234 14492 3240 14544
rect 3292 14532 3298 14544
rect 7285 14535 7343 14541
rect 7285 14532 7297 14535
rect 3292 14504 7297 14532
rect 3292 14492 3298 14504
rect 7285 14501 7297 14504
rect 7331 14501 7343 14535
rect 7285 14495 7343 14501
rect 7484 14504 7788 14532
rect 2866 14464 2872 14476
rect 2332 14436 2872 14464
rect 1670 14356 1676 14408
rect 1728 14356 1734 14408
rect 2332 14405 2360 14436
rect 2866 14424 2872 14436
rect 2924 14464 2930 14476
rect 2924 14436 3464 14464
rect 2924 14424 2930 14436
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14365 2375 14399
rect 2317 14359 2375 14365
rect 2406 14356 2412 14408
rect 2464 14396 2470 14408
rect 2501 14399 2559 14405
rect 2501 14396 2513 14399
rect 2464 14368 2513 14396
rect 2464 14356 2470 14368
rect 2501 14365 2513 14368
rect 2547 14365 2559 14399
rect 2501 14359 2559 14365
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14365 2651 14399
rect 2593 14359 2651 14365
rect 2608 14260 2636 14359
rect 3436 14328 3464 14436
rect 4062 14424 4068 14476
rect 4120 14464 4126 14476
rect 4120 14436 4384 14464
rect 4120 14424 4126 14436
rect 3970 14356 3976 14408
rect 4028 14396 4034 14408
rect 4356 14405 4384 14436
rect 4798 14424 4804 14476
rect 4856 14464 4862 14476
rect 6273 14467 6331 14473
rect 6273 14464 6285 14467
rect 4856 14436 6285 14464
rect 4856 14424 4862 14436
rect 6273 14433 6285 14436
rect 6319 14464 6331 14467
rect 7484 14464 7512 14504
rect 6319 14436 7512 14464
rect 6319 14433 6331 14436
rect 6273 14427 6331 14433
rect 7558 14424 7564 14476
rect 7616 14424 7622 14476
rect 7760 14473 7788 14504
rect 7745 14467 7803 14473
rect 7745 14433 7757 14467
rect 7791 14433 7803 14467
rect 8036 14464 8064 14572
rect 9122 14560 9128 14572
rect 9180 14560 9186 14612
rect 9309 14603 9367 14609
rect 9309 14569 9321 14603
rect 9355 14600 9367 14603
rect 9490 14600 9496 14612
rect 9355 14572 9496 14600
rect 9355 14569 9367 14572
rect 9309 14563 9367 14569
rect 9490 14560 9496 14572
rect 9548 14600 9554 14612
rect 9674 14600 9680 14612
rect 9548 14572 9680 14600
rect 9548 14560 9554 14572
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 10229 14603 10287 14609
rect 10229 14569 10241 14603
rect 10275 14600 10287 14603
rect 11514 14600 11520 14612
rect 10275 14572 11520 14600
rect 10275 14569 10287 14572
rect 10229 14563 10287 14569
rect 11514 14560 11520 14572
rect 11572 14560 11578 14612
rect 11793 14603 11851 14609
rect 11793 14569 11805 14603
rect 11839 14600 11851 14603
rect 12526 14600 12532 14612
rect 11839 14572 12532 14600
rect 11839 14569 11851 14572
rect 11793 14563 11851 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 12805 14603 12863 14609
rect 12805 14569 12817 14603
rect 12851 14600 12863 14603
rect 12986 14600 12992 14612
rect 12851 14572 12992 14600
rect 12851 14569 12863 14572
rect 12805 14563 12863 14569
rect 12986 14560 12992 14572
rect 13044 14560 13050 14612
rect 8202 14492 8208 14544
rect 8260 14532 8266 14544
rect 10873 14535 10931 14541
rect 10873 14532 10885 14535
rect 8260 14504 10885 14532
rect 8260 14492 8266 14504
rect 10873 14501 10885 14504
rect 10919 14501 10931 14535
rect 10873 14495 10931 14501
rect 10962 14492 10968 14544
rect 11020 14492 11026 14544
rect 11348 14504 12848 14532
rect 7745 14427 7803 14433
rect 7852 14436 8064 14464
rect 8665 14467 8723 14473
rect 4157 14399 4215 14405
rect 4157 14396 4169 14399
rect 4028 14368 4169 14396
rect 4028 14356 4034 14368
rect 4157 14365 4169 14368
rect 4203 14365 4215 14399
rect 4157 14359 4215 14365
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14365 4399 14399
rect 4341 14359 4399 14365
rect 4430 14356 4436 14408
rect 4488 14356 4494 14408
rect 4706 14356 4712 14408
rect 4764 14396 4770 14408
rect 4893 14399 4951 14405
rect 4764 14368 4844 14396
rect 4764 14356 4770 14368
rect 3436 14300 4752 14328
rect 4724 14272 4752 14300
rect 3973 14263 4031 14269
rect 3973 14260 3985 14263
rect 2608 14232 3985 14260
rect 3973 14229 3985 14232
rect 4019 14229 4031 14263
rect 3973 14223 4031 14229
rect 4522 14220 4528 14272
rect 4580 14220 4586 14272
rect 4706 14220 4712 14272
rect 4764 14220 4770 14272
rect 4816 14260 4844 14368
rect 4893 14365 4905 14399
rect 4939 14365 4951 14399
rect 4893 14359 4951 14365
rect 4985 14399 5043 14405
rect 4985 14365 4997 14399
rect 5031 14396 5043 14399
rect 5258 14396 5264 14408
rect 5031 14368 5264 14396
rect 5031 14365 5043 14368
rect 4985 14359 5043 14365
rect 4908 14328 4936 14359
rect 5258 14356 5264 14368
rect 5316 14396 5322 14408
rect 5994 14396 6000 14408
rect 5316 14368 6000 14396
rect 5316 14356 5322 14368
rect 5994 14356 6000 14368
rect 6052 14356 6058 14408
rect 6181 14399 6239 14405
rect 6181 14365 6193 14399
rect 6227 14365 6239 14399
rect 6181 14359 6239 14365
rect 4908 14300 5304 14328
rect 5169 14263 5227 14269
rect 5169 14260 5181 14263
rect 4816 14232 5181 14260
rect 5169 14229 5181 14232
rect 5215 14229 5227 14263
rect 5276 14260 5304 14300
rect 5810 14288 5816 14340
rect 5868 14328 5874 14340
rect 5905 14331 5963 14337
rect 5905 14328 5917 14331
rect 5868 14300 5917 14328
rect 5868 14288 5874 14300
rect 5905 14297 5917 14300
rect 5951 14297 5963 14331
rect 6196 14328 6224 14359
rect 6546 14356 6552 14408
rect 6604 14356 6610 14408
rect 6638 14356 6644 14408
rect 6696 14356 6702 14408
rect 7006 14356 7012 14408
rect 7064 14356 7070 14408
rect 7469 14399 7527 14405
rect 7469 14365 7481 14399
rect 7515 14365 7527 14399
rect 7469 14359 7527 14365
rect 6270 14328 6276 14340
rect 6196 14300 6276 14328
rect 5905 14291 5963 14297
rect 6270 14288 6276 14300
rect 6328 14288 6334 14340
rect 6822 14288 6828 14340
rect 6880 14288 6886 14340
rect 6914 14288 6920 14340
rect 6972 14288 6978 14340
rect 7484 14328 7512 14359
rect 7650 14356 7656 14408
rect 7708 14396 7714 14408
rect 7852 14396 7880 14436
rect 8665 14433 8677 14467
rect 8711 14464 8723 14467
rect 9217 14467 9275 14473
rect 8711 14436 8984 14464
rect 8711 14433 8723 14436
rect 8665 14427 8723 14433
rect 7708 14368 7880 14396
rect 7708 14356 7714 14368
rect 8294 14356 8300 14408
rect 8352 14396 8358 14408
rect 8573 14399 8631 14405
rect 8573 14396 8585 14399
rect 8352 14368 8585 14396
rect 8352 14356 8358 14368
rect 8573 14365 8585 14368
rect 8619 14365 8631 14399
rect 8573 14359 8631 14365
rect 8757 14399 8815 14405
rect 8757 14365 8769 14399
rect 8803 14365 8815 14399
rect 8757 14359 8815 14365
rect 8018 14328 8024 14340
rect 7484 14300 8024 14328
rect 8018 14288 8024 14300
rect 8076 14288 8082 14340
rect 8772 14328 8800 14359
rect 8846 14356 8852 14408
rect 8904 14396 8910 14408
rect 8956 14405 8984 14436
rect 9217 14433 9229 14467
rect 9263 14464 9275 14467
rect 10502 14464 10508 14476
rect 9263 14436 10508 14464
rect 9263 14433 9275 14436
rect 9217 14427 9275 14433
rect 8941 14399 8999 14405
rect 8941 14396 8953 14399
rect 8904 14368 8953 14396
rect 8904 14356 8910 14368
rect 8941 14365 8953 14368
rect 8987 14365 8999 14399
rect 8941 14359 8999 14365
rect 9030 14328 9036 14340
rect 8772 14300 9036 14328
rect 9030 14288 9036 14300
rect 9088 14288 9094 14340
rect 6454 14260 6460 14272
rect 5276 14232 6460 14260
rect 5169 14223 5227 14229
rect 6454 14220 6460 14232
rect 6512 14260 6518 14272
rect 9232 14260 9260 14427
rect 10502 14424 10508 14436
rect 10560 14424 10566 14476
rect 10980 14464 11008 14492
rect 10796 14436 11008 14464
rect 9398 14356 9404 14408
rect 9456 14396 9462 14408
rect 9585 14399 9643 14405
rect 9585 14396 9597 14399
rect 9456 14368 9597 14396
rect 9456 14356 9462 14368
rect 9585 14365 9597 14368
rect 9631 14365 9643 14399
rect 9585 14359 9643 14365
rect 9769 14399 9827 14405
rect 9769 14365 9781 14399
rect 9815 14365 9827 14399
rect 9769 14359 9827 14365
rect 9784 14328 9812 14359
rect 9858 14356 9864 14408
rect 9916 14356 9922 14408
rect 9950 14356 9956 14408
rect 10008 14356 10014 14408
rect 10796 14405 10824 14436
rect 10781 14399 10839 14405
rect 10781 14365 10793 14399
rect 10827 14365 10839 14399
rect 10781 14359 10839 14365
rect 10965 14399 11023 14405
rect 10965 14365 10977 14399
rect 11011 14396 11023 14399
rect 11146 14396 11152 14408
rect 11011 14368 11152 14396
rect 11011 14365 11023 14368
rect 10965 14359 11023 14365
rect 11146 14356 11152 14368
rect 11204 14356 11210 14408
rect 11348 14405 11376 14504
rect 11422 14424 11428 14476
rect 11480 14464 11486 14476
rect 11480 14436 12480 14464
rect 11480 14424 11486 14436
rect 11297 14399 11376 14405
rect 11297 14365 11309 14399
rect 11343 14368 11376 14399
rect 11633 14399 11691 14405
rect 11633 14396 11645 14399
rect 11343 14365 11355 14368
rect 11297 14359 11355 14365
rect 11629 14365 11645 14396
rect 11679 14365 11691 14399
rect 11629 14359 11691 14365
rect 9508 14300 9812 14328
rect 9508 14269 9536 14300
rect 11422 14288 11428 14340
rect 11480 14288 11486 14340
rect 11514 14288 11520 14340
rect 11572 14288 11578 14340
rect 11629 14328 11657 14359
rect 12342 14356 12348 14408
rect 12400 14356 12406 14408
rect 11624 14300 11657 14328
rect 6512 14232 9260 14260
rect 9493 14263 9551 14269
rect 6512 14220 6518 14232
rect 9493 14229 9505 14263
rect 9539 14229 9551 14263
rect 9493 14223 9551 14229
rect 10686 14220 10692 14272
rect 10744 14260 10750 14272
rect 11624 14260 11652 14300
rect 10744 14232 11652 14260
rect 12452 14260 12480 14436
rect 12710 14424 12716 14476
rect 12768 14424 12774 14476
rect 12820 14464 12848 14504
rect 12894 14492 12900 14544
rect 12952 14532 12958 14544
rect 14093 14535 14151 14541
rect 14093 14532 14105 14535
rect 12952 14504 14105 14532
rect 12952 14492 12958 14504
rect 14093 14501 14105 14504
rect 14139 14501 14151 14535
rect 15930 14532 15936 14544
rect 14093 14495 14151 14501
rect 14200 14504 15936 14532
rect 13722 14464 13728 14476
rect 12820 14436 13728 14464
rect 13722 14424 13728 14436
rect 13780 14424 13786 14476
rect 12526 14356 12532 14408
rect 12584 14356 12590 14408
rect 12621 14399 12679 14405
rect 12621 14365 12633 14399
rect 12667 14396 12679 14399
rect 12802 14396 12808 14408
rect 12667 14368 12808 14396
rect 12667 14365 12679 14368
rect 12621 14359 12679 14365
rect 12802 14356 12808 14368
rect 12860 14396 12866 14408
rect 13906 14396 13912 14408
rect 12860 14368 13912 14396
rect 12860 14356 12866 14368
rect 13906 14356 13912 14368
rect 13964 14356 13970 14408
rect 12894 14288 12900 14340
rect 12952 14288 12958 14340
rect 14200 14260 14228 14504
rect 15930 14492 15936 14504
rect 15988 14492 15994 14544
rect 16301 14535 16359 14541
rect 16301 14501 16313 14535
rect 16347 14532 16359 14535
rect 16482 14532 16488 14544
rect 16347 14504 16488 14532
rect 16347 14501 16359 14504
rect 16301 14495 16359 14501
rect 16482 14492 16488 14504
rect 16540 14492 16546 14544
rect 15562 14464 15568 14476
rect 14660 14436 15568 14464
rect 14274 14356 14280 14408
rect 14332 14356 14338 14408
rect 14660 14405 14688 14436
rect 15562 14424 15568 14436
rect 15620 14424 15626 14476
rect 15654 14424 15660 14476
rect 15712 14424 15718 14476
rect 15746 14424 15752 14476
rect 15804 14424 15810 14476
rect 16117 14467 16175 14473
rect 16117 14433 16129 14467
rect 16163 14464 16175 14467
rect 17678 14464 17684 14476
rect 16163 14436 17684 14464
rect 16163 14433 16175 14436
rect 16117 14427 16175 14433
rect 17678 14424 17684 14436
rect 17736 14424 17742 14476
rect 17770 14424 17776 14476
rect 17828 14464 17834 14476
rect 18049 14467 18107 14473
rect 18049 14464 18061 14467
rect 17828 14436 18061 14464
rect 17828 14424 17834 14436
rect 18049 14433 18061 14436
rect 18095 14433 18107 14467
rect 18049 14427 18107 14433
rect 14645 14399 14703 14405
rect 14645 14365 14657 14399
rect 14691 14365 14703 14399
rect 14645 14359 14703 14365
rect 14737 14399 14795 14405
rect 14737 14365 14749 14399
rect 14783 14396 14795 14399
rect 14826 14396 14832 14408
rect 14783 14368 14832 14396
rect 14783 14365 14795 14368
rect 14737 14359 14795 14365
rect 14826 14356 14832 14368
rect 14884 14356 14890 14408
rect 14921 14399 14979 14405
rect 14921 14365 14933 14399
rect 14967 14396 14979 14399
rect 15010 14396 15016 14408
rect 14967 14368 15016 14396
rect 14967 14365 14979 14368
rect 14921 14359 14979 14365
rect 15010 14356 15016 14368
rect 15068 14356 15074 14408
rect 15286 14356 15292 14408
rect 15344 14356 15350 14408
rect 15470 14356 15476 14408
rect 15528 14396 15534 14408
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 15528 14368 15853 14396
rect 15528 14356 15534 14368
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 15933 14399 15991 14405
rect 15933 14365 15945 14399
rect 15979 14365 15991 14399
rect 15933 14359 15991 14365
rect 14366 14288 14372 14340
rect 14424 14288 14430 14340
rect 14458 14288 14464 14340
rect 14516 14328 14522 14340
rect 15105 14331 15163 14337
rect 15105 14328 15117 14331
rect 14516 14300 15117 14328
rect 14516 14288 14522 14300
rect 15105 14297 15117 14300
rect 15151 14297 15163 14331
rect 15105 14291 15163 14297
rect 15197 14331 15255 14337
rect 15197 14297 15209 14331
rect 15243 14297 15255 14331
rect 15948 14328 15976 14359
rect 15948 14300 16528 14328
rect 15197 14291 15255 14297
rect 12452 14232 14228 14260
rect 14384 14260 14412 14288
rect 15212 14260 15240 14291
rect 14384 14232 15240 14260
rect 10744 14220 10750 14232
rect 15470 14220 15476 14272
rect 15528 14220 15534 14272
rect 16500 14260 16528 14300
rect 17310 14288 17316 14340
rect 17368 14288 17374 14340
rect 17494 14288 17500 14340
rect 17552 14328 17558 14340
rect 17773 14331 17831 14337
rect 17773 14328 17785 14331
rect 17552 14300 17785 14328
rect 17552 14288 17558 14300
rect 17773 14297 17785 14300
rect 17819 14297 17831 14331
rect 17773 14291 17831 14297
rect 17034 14260 17040 14272
rect 16500 14232 17040 14260
rect 17034 14220 17040 14232
rect 17092 14220 17098 14272
rect 1104 14170 18400 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 18400 14170
rect 1104 14096 18400 14118
rect 1578 14016 1584 14068
rect 1636 14056 1642 14068
rect 2682 14056 2688 14068
rect 1636 14028 2688 14056
rect 1636 14016 1642 14028
rect 2682 14016 2688 14028
rect 2740 14016 2746 14068
rect 4062 14016 4068 14068
rect 4120 14056 4126 14068
rect 4157 14059 4215 14065
rect 4157 14056 4169 14059
rect 4120 14028 4169 14056
rect 4120 14016 4126 14028
rect 4157 14025 4169 14028
rect 4203 14025 4215 14059
rect 4157 14019 4215 14025
rect 4430 14016 4436 14068
rect 4488 14056 4494 14068
rect 5997 14059 6055 14065
rect 5997 14056 6009 14059
rect 4488 14028 6009 14056
rect 4488 14016 4494 14028
rect 5997 14025 6009 14028
rect 6043 14025 6055 14059
rect 5997 14019 6055 14025
rect 6730 14016 6736 14068
rect 6788 14056 6794 14068
rect 8662 14056 8668 14068
rect 6788 14028 8668 14056
rect 6788 14016 6794 14028
rect 2516 13960 3188 13988
rect 1670 13880 1676 13932
rect 1728 13880 1734 13932
rect 2516 13929 2544 13960
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13889 2559 13923
rect 2501 13883 2559 13889
rect 2774 13880 2780 13932
rect 2832 13880 2838 13932
rect 3050 13880 3056 13932
rect 3108 13880 3114 13932
rect 3160 13852 3188 13960
rect 3234 13948 3240 14000
rect 3292 13948 3298 14000
rect 5074 13948 5080 14000
rect 5132 13988 5138 14000
rect 5537 13991 5595 13997
rect 5132 13960 5408 13988
rect 5132 13948 5138 13960
rect 3881 13923 3939 13929
rect 3881 13889 3893 13923
rect 3927 13920 3939 13923
rect 4522 13920 4528 13932
rect 3927 13892 4528 13920
rect 3927 13889 3939 13892
rect 3881 13883 3939 13889
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 5380 13929 5408 13960
rect 5537 13957 5549 13991
rect 5583 13988 5595 13991
rect 5626 13988 5632 14000
rect 5583 13960 5632 13988
rect 5583 13957 5595 13960
rect 5537 13951 5595 13957
rect 5626 13948 5632 13960
rect 5684 13948 5690 14000
rect 5718 13948 5724 14000
rect 5776 13997 5782 14000
rect 5776 13991 5795 13997
rect 5783 13957 5795 13991
rect 5776 13951 5795 13957
rect 5776 13948 5782 13951
rect 5169 13923 5227 13929
rect 5169 13889 5181 13923
rect 5215 13889 5227 13923
rect 5169 13883 5227 13889
rect 5261 13923 5319 13929
rect 5261 13889 5273 13923
rect 5307 13889 5319 13923
rect 5261 13883 5319 13889
rect 5353 13923 5411 13929
rect 5353 13889 5365 13923
rect 5399 13889 5411 13923
rect 5997 13923 6055 13929
rect 5997 13920 6009 13923
rect 5353 13883 5411 13889
rect 5828 13892 6009 13920
rect 4062 13852 4068 13864
rect 3160 13824 4068 13852
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 4157 13855 4215 13861
rect 4157 13821 4169 13855
rect 4203 13852 4215 13855
rect 4798 13852 4804 13864
rect 4203 13824 4804 13852
rect 4203 13821 4215 13824
rect 4157 13815 4215 13821
rect 4798 13812 4804 13824
rect 4856 13852 4862 13864
rect 5184 13852 5212 13883
rect 4856 13824 5212 13852
rect 5276 13852 5304 13883
rect 5828 13852 5856 13892
rect 5997 13889 6009 13892
rect 6043 13889 6055 13923
rect 5997 13883 6055 13889
rect 6178 13880 6184 13932
rect 6236 13880 6242 13932
rect 6914 13880 6920 13932
rect 6972 13880 6978 13932
rect 7098 13880 7104 13932
rect 7156 13880 7162 13932
rect 7392 13929 7420 14028
rect 8662 14016 8668 14028
rect 8720 14016 8726 14068
rect 9493 14059 9551 14065
rect 9493 14025 9505 14059
rect 9539 14056 9551 14059
rect 9858 14056 9864 14068
rect 9539 14028 9864 14056
rect 9539 14025 9551 14028
rect 9493 14019 9551 14025
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 11330 14016 11336 14068
rect 11388 14016 11394 14068
rect 11422 14016 11428 14068
rect 11480 14056 11486 14068
rect 11517 14059 11575 14065
rect 11517 14056 11529 14059
rect 11480 14028 11529 14056
rect 11480 14016 11486 14028
rect 11517 14025 11529 14028
rect 11563 14025 11575 14059
rect 14366 14056 14372 14068
rect 11517 14019 11575 14025
rect 14292 14028 14372 14056
rect 7650 13948 7656 14000
rect 7708 13988 7714 14000
rect 10594 13988 10600 14000
rect 7708 13960 8156 13988
rect 7708 13948 7714 13960
rect 8128 13932 8156 13960
rect 8312 13960 10600 13988
rect 7377 13923 7435 13929
rect 7377 13889 7389 13923
rect 7423 13889 7435 13923
rect 7377 13883 7435 13889
rect 7561 13923 7619 13929
rect 7561 13889 7573 13923
rect 7607 13920 7619 13923
rect 7929 13923 7987 13929
rect 7929 13920 7941 13923
rect 7607 13892 7941 13920
rect 7607 13889 7619 13892
rect 7561 13883 7619 13889
rect 7929 13889 7941 13892
rect 7975 13889 7987 13923
rect 7929 13883 7987 13889
rect 8018 13880 8024 13932
rect 8076 13880 8082 13932
rect 8110 13880 8116 13932
rect 8168 13920 8174 13932
rect 8312 13929 8340 13960
rect 10594 13948 10600 13960
rect 10652 13948 10658 14000
rect 11348 13951 11376 14016
rect 11333 13945 11391 13951
rect 8205 13923 8263 13929
rect 8205 13920 8217 13923
rect 8168 13892 8217 13920
rect 8168 13880 8174 13892
rect 8205 13889 8217 13892
rect 8251 13889 8263 13923
rect 8205 13883 8263 13889
rect 8297 13923 8355 13929
rect 8297 13889 8309 13923
rect 8343 13889 8355 13923
rect 8297 13883 8355 13889
rect 8570 13880 8576 13932
rect 8628 13880 8634 13932
rect 8846 13880 8852 13932
rect 8904 13880 8910 13932
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13889 8999 13923
rect 8941 13883 8999 13889
rect 6546 13852 6552 13864
rect 5276 13824 5856 13852
rect 4856 13812 4862 13824
rect 1486 13676 1492 13728
rect 1544 13676 1550 13728
rect 2314 13676 2320 13728
rect 2372 13676 2378 13728
rect 2866 13676 2872 13728
rect 2924 13676 2930 13728
rect 3970 13676 3976 13728
rect 4028 13676 4034 13728
rect 5718 13725 5724 13728
rect 5712 13716 5724 13725
rect 5679 13688 5724 13716
rect 5712 13679 5724 13688
rect 5718 13676 5724 13679
rect 5776 13676 5782 13728
rect 5828 13716 5856 13824
rect 5920 13824 6552 13852
rect 5920 13793 5948 13824
rect 6546 13812 6552 13824
rect 6604 13852 6610 13864
rect 7193 13855 7251 13861
rect 7193 13852 7205 13855
rect 6604 13824 7205 13852
rect 6604 13812 6610 13824
rect 7193 13821 7205 13824
rect 7239 13821 7251 13855
rect 7193 13815 7251 13821
rect 7285 13855 7343 13861
rect 7285 13821 7297 13855
rect 7331 13852 7343 13855
rect 7834 13852 7840 13864
rect 7331 13824 7840 13852
rect 7331 13821 7343 13824
rect 7285 13815 7343 13821
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 8956 13852 8984 13883
rect 9398 13880 9404 13932
rect 9456 13880 9462 13932
rect 9582 13880 9588 13932
rect 9640 13880 9646 13932
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 10045 13923 10103 13929
rect 10045 13920 10057 13923
rect 9916 13892 10057 13920
rect 9916 13880 9922 13892
rect 10045 13889 10057 13892
rect 10091 13920 10103 13923
rect 10778 13920 10784 13932
rect 10091 13892 10784 13920
rect 10091 13889 10103 13892
rect 10045 13883 10103 13889
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 11057 13923 11115 13929
rect 11057 13889 11069 13923
rect 11103 13889 11115 13923
rect 11057 13883 11115 13889
rect 11241 13923 11299 13929
rect 11241 13889 11253 13923
rect 11287 13889 11299 13923
rect 11333 13911 11345 13945
rect 11379 13911 11391 13945
rect 11333 13905 11391 13911
rect 11241 13883 11299 13889
rect 8312 13824 8984 13852
rect 5905 13787 5963 13793
rect 5905 13753 5917 13787
rect 5951 13753 5963 13787
rect 5905 13747 5963 13753
rect 7650 13716 7656 13728
rect 5828 13688 7656 13716
rect 7650 13676 7656 13688
rect 7708 13716 7714 13728
rect 8312 13716 8340 13824
rect 8478 13744 8484 13796
rect 8536 13744 8542 13796
rect 8570 13744 8576 13796
rect 8628 13784 8634 13796
rect 11072 13784 11100 13883
rect 11256 13852 11284 13883
rect 11698 13880 11704 13932
rect 11756 13880 11762 13932
rect 11793 13923 11851 13929
rect 11793 13889 11805 13923
rect 11839 13920 11851 13923
rect 13078 13920 13084 13932
rect 11839 13892 13084 13920
rect 11839 13889 11851 13892
rect 11793 13883 11851 13889
rect 11808 13852 11836 13883
rect 13078 13880 13084 13892
rect 13136 13920 13142 13932
rect 13354 13920 13360 13932
rect 13136 13892 13360 13920
rect 13136 13880 13142 13892
rect 13354 13880 13360 13892
rect 13412 13880 13418 13932
rect 13446 13880 13452 13932
rect 13504 13920 13510 13932
rect 14292 13929 14320 14028
rect 14366 14016 14372 14028
rect 14424 14016 14430 14068
rect 14737 14059 14795 14065
rect 14737 14025 14749 14059
rect 14783 14056 14795 14059
rect 16758 14056 16764 14068
rect 14783 14028 16764 14056
rect 14783 14025 14795 14028
rect 14737 14019 14795 14025
rect 16758 14016 16764 14028
rect 16816 14016 16822 14068
rect 16942 14016 16948 14068
rect 17000 14016 17006 14068
rect 17034 14016 17040 14068
rect 17092 14016 17098 14068
rect 17494 14016 17500 14068
rect 17552 14016 17558 14068
rect 17954 14016 17960 14068
rect 18012 14016 18018 14068
rect 14826 13988 14832 14000
rect 14476 13960 14832 13988
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 13504 13892 14289 13920
rect 13504 13880 13510 13892
rect 14277 13889 14289 13892
rect 14323 13889 14335 13923
rect 14277 13883 14335 13889
rect 14366 13880 14372 13932
rect 14424 13880 14430 13932
rect 11256 13824 11836 13852
rect 12158 13812 12164 13864
rect 12216 13812 12222 13864
rect 14093 13855 14151 13861
rect 14093 13821 14105 13855
rect 14139 13821 14151 13855
rect 14093 13815 14151 13821
rect 11974 13784 11980 13796
rect 8628 13756 11008 13784
rect 11072 13756 11980 13784
rect 8628 13744 8634 13756
rect 7708 13688 8340 13716
rect 8665 13719 8723 13725
rect 7708 13676 7714 13688
rect 8665 13685 8677 13719
rect 8711 13716 8723 13719
rect 8754 13716 8760 13728
rect 8711 13688 8760 13716
rect 8711 13685 8723 13688
rect 8665 13679 8723 13685
rect 8754 13676 8760 13688
rect 8812 13716 8818 13728
rect 9030 13716 9036 13728
rect 8812 13688 9036 13716
rect 8812 13676 8818 13688
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 9125 13719 9183 13725
rect 9125 13685 9137 13719
rect 9171 13716 9183 13719
rect 9214 13716 9220 13728
rect 9171 13688 9220 13716
rect 9171 13685 9183 13688
rect 9125 13679 9183 13685
rect 9214 13676 9220 13688
rect 9272 13676 9278 13728
rect 9766 13676 9772 13728
rect 9824 13676 9830 13728
rect 10686 13676 10692 13728
rect 10744 13716 10750 13728
rect 10873 13719 10931 13725
rect 10873 13716 10885 13719
rect 10744 13688 10885 13716
rect 10744 13676 10750 13688
rect 10873 13685 10885 13688
rect 10919 13685 10931 13719
rect 10980 13716 11008 13756
rect 11974 13744 11980 13756
rect 12032 13744 12038 13796
rect 14108 13784 14136 13815
rect 14182 13812 14188 13864
rect 14240 13812 14246 13864
rect 14476 13784 14504 13960
rect 14826 13948 14832 13960
rect 14884 13948 14890 14000
rect 15470 13948 15476 14000
rect 15528 13988 15534 14000
rect 15528 13960 17264 13988
rect 15528 13948 15534 13960
rect 14642 13880 14648 13932
rect 14700 13880 14706 13932
rect 14918 13880 14924 13932
rect 14976 13880 14982 13932
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13920 15071 13923
rect 15378 13920 15384 13932
rect 15059 13892 15384 13920
rect 15059 13889 15071 13892
rect 15013 13883 15071 13889
rect 15378 13880 15384 13892
rect 15436 13880 15442 13932
rect 16209 13923 16267 13929
rect 15580 13892 16160 13920
rect 14553 13855 14611 13861
rect 14553 13821 14565 13855
rect 14599 13852 14611 13855
rect 14599 13824 14780 13852
rect 14599 13821 14611 13824
rect 14553 13815 14611 13821
rect 14108 13756 14504 13784
rect 14752 13784 14780 13824
rect 14826 13812 14832 13864
rect 14884 13812 14890 13864
rect 15580 13852 15608 13892
rect 14936 13824 15608 13852
rect 14936 13784 14964 13824
rect 15654 13812 15660 13864
rect 15712 13812 15718 13864
rect 15933 13855 15991 13861
rect 15933 13821 15945 13855
rect 15979 13852 15991 13855
rect 16022 13852 16028 13864
rect 15979 13824 16028 13852
rect 15979 13821 15991 13824
rect 15933 13815 15991 13821
rect 16022 13812 16028 13824
rect 16080 13812 16086 13864
rect 16132 13852 16160 13892
rect 16209 13889 16221 13923
rect 16255 13920 16267 13923
rect 16574 13920 16580 13932
rect 16255 13892 16580 13920
rect 16255 13889 16267 13892
rect 16209 13883 16267 13889
rect 16574 13880 16580 13892
rect 16632 13880 16638 13932
rect 17236 13929 17264 13960
rect 16669 13923 16727 13929
rect 16669 13889 16681 13923
rect 16715 13889 16727 13923
rect 17037 13923 17095 13929
rect 17037 13920 17049 13923
rect 16669 13883 16727 13889
rect 16960 13892 17049 13920
rect 16684 13852 16712 13883
rect 16132 13824 16712 13852
rect 16758 13812 16764 13864
rect 16816 13852 16822 13864
rect 16960 13861 16988 13892
rect 17037 13889 17049 13892
rect 17083 13889 17095 13923
rect 17037 13883 17095 13889
rect 17221 13923 17279 13929
rect 17221 13889 17233 13923
rect 17267 13889 17279 13923
rect 17221 13883 17279 13889
rect 17313 13923 17371 13929
rect 17313 13889 17325 13923
rect 17359 13920 17371 13923
rect 17402 13920 17408 13932
rect 17359 13892 17408 13920
rect 17359 13889 17371 13892
rect 17313 13883 17371 13889
rect 17402 13880 17408 13892
rect 17460 13880 17466 13932
rect 17497 13923 17555 13929
rect 17497 13889 17509 13923
rect 17543 13920 17555 13923
rect 17586 13920 17592 13932
rect 17543 13892 17592 13920
rect 17543 13889 17555 13892
rect 17497 13883 17555 13889
rect 17586 13880 17592 13892
rect 17644 13880 17650 13932
rect 17678 13880 17684 13932
rect 17736 13920 17742 13932
rect 17773 13923 17831 13929
rect 17773 13920 17785 13923
rect 17736 13892 17785 13920
rect 17736 13880 17742 13892
rect 17773 13889 17785 13892
rect 17819 13889 17831 13923
rect 17773 13883 17831 13889
rect 16945 13855 17003 13861
rect 16945 13852 16957 13855
rect 16816 13824 16957 13852
rect 16816 13812 16822 13824
rect 16945 13821 16957 13824
rect 16991 13821 17003 13855
rect 16945 13815 17003 13821
rect 14752 13756 14964 13784
rect 15102 13744 15108 13796
rect 15160 13784 15166 13796
rect 15160 13756 16804 13784
rect 15160 13744 15166 13756
rect 11514 13716 11520 13728
rect 10980 13688 11520 13716
rect 10873 13679 10931 13685
rect 11514 13676 11520 13688
rect 11572 13676 11578 13728
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 14826 13716 14832 13728
rect 12768 13688 14832 13716
rect 12768 13676 12774 13688
rect 14826 13676 14832 13688
rect 14884 13676 14890 13728
rect 16776 13725 16804 13756
rect 16761 13719 16819 13725
rect 16761 13685 16773 13719
rect 16807 13685 16819 13719
rect 16761 13679 16819 13685
rect 1104 13626 18400 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 18400 13626
rect 1104 13552 18400 13574
rect 2866 13512 2872 13524
rect 1504 13484 2872 13512
rect 1504 13317 1532 13484
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 3326 13472 3332 13524
rect 3384 13472 3390 13524
rect 3878 13472 3884 13524
rect 3936 13512 3942 13524
rect 4157 13515 4215 13521
rect 4157 13512 4169 13515
rect 3936 13484 4169 13512
rect 3936 13472 3942 13484
rect 4157 13481 4169 13484
rect 4203 13512 4215 13515
rect 4890 13512 4896 13524
rect 4203 13484 4896 13512
rect 4203 13481 4215 13484
rect 4157 13475 4215 13481
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 5442 13472 5448 13524
rect 5500 13512 5506 13524
rect 6454 13512 6460 13524
rect 5500 13484 6460 13512
rect 5500 13472 5506 13484
rect 6454 13472 6460 13484
rect 6512 13472 6518 13524
rect 7098 13472 7104 13524
rect 7156 13472 7162 13524
rect 7190 13472 7196 13524
rect 7248 13512 7254 13524
rect 7285 13515 7343 13521
rect 7285 13512 7297 13515
rect 7248 13484 7297 13512
rect 7248 13472 7254 13484
rect 7285 13481 7297 13484
rect 7331 13481 7343 13515
rect 7285 13475 7343 13481
rect 8018 13472 8024 13524
rect 8076 13512 8082 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 8076 13484 8953 13512
rect 8076 13472 8082 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 10686 13512 10692 13524
rect 8941 13475 8999 13481
rect 9048 13484 10692 13512
rect 1765 13447 1823 13453
rect 1765 13413 1777 13447
rect 1811 13444 1823 13447
rect 2593 13447 2651 13453
rect 1811 13416 2544 13444
rect 1811 13413 1823 13416
rect 1765 13407 1823 13413
rect 2041 13379 2099 13385
rect 2041 13345 2053 13379
rect 2087 13376 2099 13379
rect 2314 13376 2320 13388
rect 2087 13348 2320 13376
rect 2087 13345 2099 13348
rect 2041 13339 2099 13345
rect 2314 13336 2320 13348
rect 2372 13336 2378 13388
rect 2516 13376 2544 13416
rect 2593 13413 2605 13447
rect 2639 13444 2651 13447
rect 3344 13444 3372 13472
rect 2639 13416 3372 13444
rect 8665 13447 8723 13453
rect 2639 13413 2651 13416
rect 2593 13407 2651 13413
rect 8665 13413 8677 13447
rect 8711 13444 8723 13447
rect 8846 13444 8852 13456
rect 8711 13416 8852 13444
rect 8711 13413 8723 13416
rect 8665 13407 8723 13413
rect 8846 13404 8852 13416
rect 8904 13404 8910 13456
rect 2516 13348 3004 13376
rect 1489 13311 1547 13317
rect 1489 13277 1501 13311
rect 1535 13277 1547 13311
rect 1489 13271 1547 13277
rect 1578 13268 1584 13320
rect 1636 13268 1642 13320
rect 1765 13311 1823 13317
rect 1765 13277 1777 13311
rect 1811 13308 1823 13311
rect 2498 13308 2504 13320
rect 1811 13280 2504 13308
rect 1811 13277 1823 13280
rect 1765 13271 1823 13277
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 2866 13308 2872 13320
rect 2608 13280 2872 13308
rect 2608 13249 2636 13280
rect 2866 13268 2872 13280
rect 2924 13268 2930 13320
rect 2976 13317 3004 13348
rect 3050 13336 3056 13388
rect 3108 13376 3114 13388
rect 3602 13376 3608 13388
rect 3108 13348 3608 13376
rect 3108 13336 3114 13348
rect 3602 13336 3608 13348
rect 3660 13376 3666 13388
rect 6914 13376 6920 13388
rect 3660 13348 4016 13376
rect 3660 13336 3666 13348
rect 2964 13311 3022 13317
rect 2964 13277 2976 13311
rect 3010 13277 3022 13311
rect 2964 13271 3022 13277
rect 3142 13268 3148 13320
rect 3200 13268 3206 13320
rect 3786 13268 3792 13320
rect 3844 13268 3850 13320
rect 3988 13317 4016 13348
rect 5276 13348 6920 13376
rect 5276 13317 5304 13348
rect 6914 13336 6920 13348
rect 6972 13336 6978 13388
rect 9048 13376 9076 13484
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 10781 13515 10839 13521
rect 10781 13481 10793 13515
rect 10827 13512 10839 13515
rect 10870 13512 10876 13524
rect 10827 13484 10876 13512
rect 10827 13481 10839 13484
rect 10781 13475 10839 13481
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 13173 13515 13231 13521
rect 13173 13512 13185 13515
rect 11204 13484 13185 13512
rect 11204 13472 11210 13484
rect 13173 13481 13185 13484
rect 13219 13481 13231 13515
rect 13173 13475 13231 13481
rect 9214 13444 9220 13456
rect 9140 13416 9220 13444
rect 9140 13385 9168 13416
rect 9214 13404 9220 13416
rect 9272 13404 9278 13456
rect 10042 13404 10048 13456
rect 10100 13444 10106 13456
rect 10962 13444 10968 13456
rect 10100 13416 10968 13444
rect 10100 13404 10106 13416
rect 10962 13404 10968 13416
rect 11020 13444 11026 13456
rect 12805 13447 12863 13453
rect 11020 13416 11284 13444
rect 11020 13404 11026 13416
rect 7668 13348 9076 13376
rect 9125 13379 9183 13385
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13277 4031 13311
rect 3973 13271 4031 13277
rect 5261 13311 5319 13317
rect 5261 13277 5273 13311
rect 5307 13277 5319 13311
rect 5261 13271 5319 13277
rect 5445 13311 5503 13317
rect 5445 13277 5457 13311
rect 5491 13308 5503 13311
rect 6362 13308 6368 13320
rect 5491 13280 6368 13308
rect 5491 13277 5503 13280
rect 5445 13271 5503 13277
rect 6362 13268 6368 13280
rect 6420 13268 6426 13320
rect 7668 13317 7696 13348
rect 9125 13345 9137 13379
rect 9171 13345 9183 13379
rect 9125 13339 9183 13345
rect 9306 13336 9312 13388
rect 9364 13376 9370 13388
rect 11256 13385 11284 13416
rect 12805 13413 12817 13447
rect 12851 13444 12863 13447
rect 12894 13444 12900 13456
rect 12851 13416 12900 13444
rect 12851 13413 12863 13416
rect 12805 13407 12863 13413
rect 12894 13404 12900 13416
rect 12952 13404 12958 13456
rect 13188 13444 13216 13475
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 15381 13515 15439 13521
rect 15381 13512 15393 13515
rect 15344 13484 15393 13512
rect 15344 13472 15350 13484
rect 15381 13481 15393 13484
rect 15427 13481 15439 13515
rect 15381 13475 15439 13481
rect 16025 13515 16083 13521
rect 16025 13481 16037 13515
rect 16071 13512 16083 13515
rect 16114 13512 16120 13524
rect 16071 13484 16120 13512
rect 16071 13481 16083 13484
rect 16025 13475 16083 13481
rect 16114 13472 16120 13484
rect 16172 13472 16178 13524
rect 17770 13472 17776 13524
rect 17828 13472 17834 13524
rect 13188 13416 13584 13444
rect 9585 13379 9643 13385
rect 9585 13376 9597 13379
rect 9364 13348 9597 13376
rect 9364 13336 9370 13348
rect 9585 13345 9597 13348
rect 9631 13345 9643 13379
rect 9585 13339 9643 13345
rect 9677 13379 9735 13385
rect 9677 13345 9689 13379
rect 9723 13345 9735 13379
rect 9677 13339 9735 13345
rect 9861 13379 9919 13385
rect 9861 13345 9873 13379
rect 9907 13376 9919 13379
rect 10505 13379 10563 13385
rect 10505 13376 10517 13379
rect 9907 13348 10517 13376
rect 9907 13345 9919 13348
rect 9861 13339 9919 13345
rect 10505 13345 10517 13348
rect 10551 13376 10563 13379
rect 11149 13379 11207 13385
rect 11149 13376 11161 13379
rect 10551 13348 11161 13376
rect 10551 13345 10563 13348
rect 10505 13339 10563 13345
rect 11149 13345 11161 13348
rect 11195 13345 11207 13379
rect 11149 13339 11207 13345
rect 11241 13379 11299 13385
rect 11241 13345 11253 13379
rect 11287 13376 11299 13379
rect 13078 13376 13084 13388
rect 11287 13348 13084 13376
rect 11287 13345 11299 13348
rect 11241 13339 11299 13345
rect 7377 13311 7435 13317
rect 7377 13277 7389 13311
rect 7423 13277 7435 13311
rect 7377 13271 7435 13277
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13277 7711 13311
rect 7653 13271 7711 13277
rect 2593 13243 2651 13249
rect 2593 13209 2605 13243
rect 2639 13209 2651 13243
rect 3421 13243 3479 13249
rect 3421 13240 3433 13243
rect 2593 13203 2651 13209
rect 2700 13212 3433 13240
rect 1857 13175 1915 13181
rect 1857 13141 1869 13175
rect 1903 13172 1915 13175
rect 1946 13172 1952 13184
rect 1903 13144 1952 13172
rect 1903 13141 1915 13144
rect 1857 13135 1915 13141
rect 1946 13132 1952 13144
rect 2004 13132 2010 13184
rect 2133 13175 2191 13181
rect 2133 13141 2145 13175
rect 2179 13172 2191 13175
rect 2700 13172 2728 13212
rect 3421 13209 3433 13212
rect 3467 13240 3479 13243
rect 5353 13243 5411 13249
rect 5353 13240 5365 13243
rect 3467 13212 5365 13240
rect 3467 13209 3479 13212
rect 3421 13203 3479 13209
rect 5353 13209 5365 13212
rect 5399 13209 5411 13243
rect 5810 13240 5816 13252
rect 5353 13203 5411 13209
rect 5460 13212 5816 13240
rect 2179 13144 2728 13172
rect 2777 13175 2835 13181
rect 2179 13141 2191 13144
rect 2133 13135 2191 13141
rect 2777 13141 2789 13175
rect 2823 13172 2835 13175
rect 2866 13172 2872 13184
rect 2823 13144 2872 13172
rect 2823 13141 2835 13144
rect 2777 13135 2835 13141
rect 2866 13132 2872 13144
rect 2924 13132 2930 13184
rect 4246 13132 4252 13184
rect 4304 13172 4310 13184
rect 5460 13172 5488 13212
rect 5810 13200 5816 13212
rect 5868 13240 5874 13252
rect 7006 13240 7012 13252
rect 5868 13212 7012 13240
rect 5868 13200 5874 13212
rect 7006 13200 7012 13212
rect 7064 13200 7070 13252
rect 7392 13240 7420 13271
rect 8570 13268 8576 13320
rect 8628 13268 8634 13320
rect 8757 13311 8815 13317
rect 8757 13277 8769 13311
rect 8803 13277 8815 13311
rect 8757 13271 8815 13277
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13308 9275 13311
rect 9692 13308 9720 13339
rect 13078 13336 13084 13348
rect 13136 13336 13142 13388
rect 13556 13376 13584 13416
rect 15010 13404 15016 13456
rect 15068 13444 15074 13456
rect 17402 13444 17408 13456
rect 15068 13416 17408 13444
rect 15068 13404 15074 13416
rect 17402 13404 17408 13416
rect 17460 13404 17466 13456
rect 15746 13376 15752 13388
rect 13188 13348 13400 13376
rect 9263 13280 9720 13308
rect 9953 13311 10011 13317
rect 9263 13277 9275 13280
rect 9217 13271 9275 13277
rect 9953 13277 9965 13311
rect 9999 13277 10011 13311
rect 9953 13271 10011 13277
rect 7926 13240 7932 13252
rect 7392 13212 7932 13240
rect 7926 13200 7932 13212
rect 7984 13200 7990 13252
rect 4304 13144 5488 13172
rect 4304 13132 4310 13144
rect 6822 13132 6828 13184
rect 6880 13172 6886 13184
rect 8570 13172 8576 13184
rect 6880 13144 8576 13172
rect 6880 13132 6886 13144
rect 8570 13132 8576 13144
rect 8628 13132 8634 13184
rect 8772 13172 8800 13271
rect 8846 13200 8852 13252
rect 8904 13240 8910 13252
rect 9306 13240 9312 13252
rect 8904 13212 9312 13240
rect 8904 13200 8910 13212
rect 9306 13200 9312 13212
rect 9364 13200 9370 13252
rect 9490 13200 9496 13252
rect 9548 13200 9554 13252
rect 9582 13200 9588 13252
rect 9640 13240 9646 13252
rect 9968 13240 9996 13271
rect 10042 13268 10048 13320
rect 10100 13268 10106 13320
rect 10137 13311 10195 13317
rect 10137 13277 10149 13311
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 9640 13212 9996 13240
rect 9640 13200 9646 13212
rect 9674 13172 9680 13184
rect 8772 13144 9680 13172
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 10152 13172 10180 13271
rect 10410 13268 10416 13320
rect 10468 13268 10474 13320
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13277 10655 13311
rect 10597 13271 10655 13277
rect 9824 13144 10180 13172
rect 10612 13172 10640 13271
rect 10686 13268 10692 13320
rect 10744 13308 10750 13320
rect 10965 13311 11023 13317
rect 10965 13308 10977 13311
rect 10744 13280 10977 13308
rect 10744 13268 10750 13280
rect 10965 13277 10977 13280
rect 11011 13277 11023 13311
rect 10965 13271 11023 13277
rect 11057 13311 11115 13317
rect 11057 13277 11069 13311
rect 11103 13277 11115 13311
rect 11057 13271 11115 13277
rect 11073 13240 11101 13271
rect 12986 13268 12992 13320
rect 13044 13308 13050 13320
rect 13188 13308 13216 13348
rect 13372 13317 13400 13348
rect 13556 13348 15752 13376
rect 13556 13317 13584 13348
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 13044 13280 13216 13308
rect 13265 13311 13323 13317
rect 13044 13268 13050 13280
rect 13265 13277 13277 13311
rect 13311 13277 13323 13311
rect 13265 13271 13323 13277
rect 13357 13311 13415 13317
rect 13357 13277 13369 13311
rect 13403 13277 13415 13311
rect 13357 13271 13415 13277
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13277 13599 13311
rect 13541 13271 13599 13277
rect 12250 13240 12256 13252
rect 11073 13212 12256 13240
rect 12250 13200 12256 13212
rect 12308 13200 12314 13252
rect 12710 13172 12716 13184
rect 10612 13144 12716 13172
rect 9824 13132 9830 13144
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 13280 13172 13308 13271
rect 13814 13268 13820 13320
rect 13872 13308 13878 13320
rect 14734 13308 14740 13320
rect 13872 13280 14740 13308
rect 13872 13268 13878 13280
rect 14734 13268 14740 13280
rect 14792 13308 14798 13320
rect 14921 13311 14979 13317
rect 14921 13308 14933 13311
rect 14792 13280 14933 13308
rect 14792 13268 14798 13280
rect 14921 13277 14933 13280
rect 14967 13308 14979 13311
rect 15010 13308 15016 13320
rect 14967 13280 15016 13308
rect 14967 13277 14979 13280
rect 14921 13271 14979 13277
rect 15010 13268 15016 13280
rect 15068 13268 15074 13320
rect 15197 13311 15255 13317
rect 15197 13277 15209 13311
rect 15243 13308 15255 13311
rect 15654 13308 15660 13320
rect 15243 13280 15660 13308
rect 15243 13277 15255 13280
rect 15197 13271 15255 13277
rect 14274 13200 14280 13252
rect 14332 13240 14338 13252
rect 15212 13240 15240 13271
rect 15654 13268 15660 13280
rect 15712 13268 15718 13320
rect 15841 13311 15899 13317
rect 15841 13277 15853 13311
rect 15887 13308 15899 13311
rect 15930 13308 15936 13320
rect 15887 13280 15936 13308
rect 15887 13277 15899 13280
rect 15841 13271 15899 13277
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 14332 13212 15240 13240
rect 14332 13200 14338 13212
rect 15286 13200 15292 13252
rect 15344 13240 15350 13252
rect 16301 13243 16359 13249
rect 16301 13240 16313 13243
rect 15344 13212 16313 13240
rect 15344 13200 15350 13212
rect 16301 13209 16313 13212
rect 16347 13209 16359 13243
rect 16301 13203 16359 13209
rect 13354 13172 13360 13184
rect 13280 13144 13360 13172
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 13541 13175 13599 13181
rect 13541 13141 13553 13175
rect 13587 13172 13599 13175
rect 13722 13172 13728 13184
rect 13587 13144 13728 13172
rect 13587 13141 13599 13144
rect 13541 13135 13599 13141
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 15010 13132 15016 13184
rect 15068 13132 15074 13184
rect 15654 13132 15660 13184
rect 15712 13172 15718 13184
rect 16390 13172 16396 13184
rect 15712 13144 16396 13172
rect 15712 13132 15718 13144
rect 16390 13132 16396 13144
rect 16448 13132 16454 13184
rect 1104 13082 18400 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 18400 13082
rect 1104 13008 18400 13030
rect 1489 12971 1547 12977
rect 1489 12937 1501 12971
rect 1535 12968 1547 12971
rect 1670 12968 1676 12980
rect 1535 12940 1676 12968
rect 1535 12937 1547 12940
rect 1489 12931 1547 12937
rect 1670 12928 1676 12940
rect 1728 12928 1734 12980
rect 1946 12928 1952 12980
rect 2004 12928 2010 12980
rect 2593 12971 2651 12977
rect 2593 12937 2605 12971
rect 2639 12968 2651 12971
rect 2682 12968 2688 12980
rect 2639 12940 2688 12968
rect 2639 12937 2651 12940
rect 2593 12931 2651 12937
rect 2682 12928 2688 12940
rect 2740 12928 2746 12980
rect 3326 12928 3332 12980
rect 3384 12968 3390 12980
rect 3605 12971 3663 12977
rect 3605 12968 3617 12971
rect 3384 12940 3617 12968
rect 3384 12928 3390 12940
rect 3605 12937 3617 12940
rect 3651 12937 3663 12971
rect 5534 12968 5540 12980
rect 3605 12931 3663 12937
rect 4540 12940 5540 12968
rect 1857 12903 1915 12909
rect 1857 12869 1869 12903
rect 1903 12900 1915 12903
rect 2866 12900 2872 12912
rect 1903 12872 2872 12900
rect 1903 12869 1915 12872
rect 1857 12863 1915 12869
rect 2866 12860 2872 12872
rect 2924 12860 2930 12912
rect 2961 12903 3019 12909
rect 2961 12869 2973 12903
rect 3007 12900 3019 12903
rect 3510 12900 3516 12912
rect 3007 12872 3516 12900
rect 3007 12869 3019 12872
rect 2961 12863 3019 12869
rect 3344 12844 3372 12872
rect 3510 12860 3516 12872
rect 3568 12860 3574 12912
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12801 2835 12835
rect 2777 12795 2835 12801
rect 2038 12724 2044 12776
rect 2096 12764 2102 12776
rect 2406 12764 2412 12776
rect 2096 12736 2412 12764
rect 2096 12724 2102 12736
rect 2406 12724 2412 12736
rect 2464 12724 2470 12776
rect 2792 12764 2820 12795
rect 3050 12792 3056 12844
rect 3108 12792 3114 12844
rect 3326 12792 3332 12844
rect 3384 12792 3390 12844
rect 3789 12835 3847 12841
rect 3789 12801 3801 12835
rect 3835 12801 3847 12835
rect 3789 12795 3847 12801
rect 3142 12764 3148 12776
rect 2792 12736 3148 12764
rect 3142 12724 3148 12736
rect 3200 12724 3206 12776
rect 3234 12724 3240 12776
rect 3292 12764 3298 12776
rect 3804 12764 3832 12795
rect 3878 12792 3884 12844
rect 3936 12792 3942 12844
rect 4065 12835 4123 12841
rect 4065 12801 4077 12835
rect 4111 12832 4123 12835
rect 4154 12832 4160 12844
rect 4111 12804 4160 12832
rect 4111 12801 4123 12804
rect 4065 12795 4123 12801
rect 4154 12792 4160 12804
rect 4212 12792 4218 12844
rect 4246 12792 4252 12844
rect 4304 12792 4310 12844
rect 4540 12832 4568 12940
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 6362 12928 6368 12980
rect 6420 12928 6426 12980
rect 8864 12940 12020 12968
rect 4614 12860 4620 12912
rect 4672 12900 4678 12912
rect 5721 12903 5779 12909
rect 4672 12872 4936 12900
rect 4672 12860 4678 12872
rect 4908 12844 4936 12872
rect 5721 12869 5733 12903
rect 5767 12900 5779 12903
rect 6851 12903 6909 12909
rect 6851 12900 6863 12903
rect 5767 12872 6863 12900
rect 5767 12869 5779 12872
rect 5721 12863 5779 12869
rect 6851 12869 6863 12872
rect 6897 12869 6909 12903
rect 6851 12863 6909 12869
rect 4709 12835 4767 12841
rect 4709 12832 4721 12835
rect 4540 12804 4721 12832
rect 4709 12801 4721 12804
rect 4755 12801 4767 12835
rect 4709 12795 4767 12801
rect 4890 12792 4896 12844
rect 4948 12792 4954 12844
rect 5074 12792 5080 12844
rect 5132 12792 5138 12844
rect 5902 12792 5908 12844
rect 5960 12792 5966 12844
rect 6086 12792 6092 12844
rect 6144 12792 6150 12844
rect 6454 12792 6460 12844
rect 6512 12832 6518 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6512 12804 6561 12832
rect 6512 12792 6518 12804
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12801 6699 12835
rect 6641 12795 6699 12801
rect 3292 12736 3832 12764
rect 3973 12767 4031 12773
rect 3292 12724 3298 12736
rect 3973 12733 3985 12767
rect 4019 12764 4031 12767
rect 4985 12767 5043 12773
rect 4985 12764 4997 12767
rect 4019 12736 4997 12764
rect 4019 12733 4031 12736
rect 3973 12727 4031 12733
rect 4985 12733 4997 12736
rect 5031 12733 5043 12767
rect 4985 12727 5043 12733
rect 6178 12724 6184 12776
rect 6236 12724 6242 12776
rect 6656 12764 6684 12795
rect 6730 12792 6736 12844
rect 6788 12792 6794 12844
rect 7009 12835 7067 12841
rect 7009 12801 7021 12835
rect 7055 12832 7067 12835
rect 8864 12832 8892 12940
rect 9033 12903 9091 12909
rect 9033 12869 9045 12903
rect 9079 12900 9091 12903
rect 9214 12900 9220 12912
rect 9079 12872 9220 12900
rect 9079 12869 9091 12872
rect 9033 12863 9091 12869
rect 9214 12860 9220 12872
rect 9272 12900 9278 12912
rect 9582 12900 9588 12912
rect 9272 12872 9588 12900
rect 9272 12860 9278 12872
rect 9582 12860 9588 12872
rect 9640 12860 9646 12912
rect 9674 12860 9680 12912
rect 9732 12900 9738 12912
rect 10410 12900 10416 12912
rect 9732 12872 10416 12900
rect 9732 12860 9738 12872
rect 7055 12804 8892 12832
rect 8941 12835 8999 12841
rect 7055 12801 7067 12804
rect 7009 12795 7067 12801
rect 8941 12801 8953 12835
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 6914 12764 6920 12776
rect 6656 12736 6920 12764
rect 6914 12724 6920 12736
rect 6972 12724 6978 12776
rect 7098 12724 7104 12776
rect 7156 12764 7162 12776
rect 8956 12764 8984 12795
rect 9122 12792 9128 12844
rect 9180 12832 9186 12844
rect 9306 12832 9312 12844
rect 9180 12804 9312 12832
rect 9180 12792 9186 12804
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 9784 12841 9812 12872
rect 10410 12860 10416 12872
rect 10468 12860 10474 12912
rect 10594 12860 10600 12912
rect 10652 12900 10658 12912
rect 11517 12903 11575 12909
rect 11517 12900 11529 12903
rect 10652 12872 11529 12900
rect 10652 12860 10658 12872
rect 11517 12869 11529 12872
rect 11563 12869 11575 12903
rect 11992 12900 12020 12940
rect 12342 12928 12348 12980
rect 12400 12968 12406 12980
rect 12986 12968 12992 12980
rect 12400 12940 12992 12968
rect 12400 12928 12406 12940
rect 12986 12928 12992 12940
rect 13044 12928 13050 12980
rect 15933 12971 15991 12977
rect 15933 12937 15945 12971
rect 15979 12937 15991 12971
rect 15933 12931 15991 12937
rect 11992 12872 13860 12900
rect 11517 12863 11575 12869
rect 9769 12835 9827 12841
rect 9769 12801 9781 12835
rect 9815 12801 9827 12835
rect 9769 12795 9827 12801
rect 9861 12835 9919 12841
rect 9861 12801 9873 12835
rect 9907 12832 9919 12835
rect 9907 12804 10640 12832
rect 9907 12801 9919 12804
rect 9861 12795 9919 12801
rect 7156 12736 8984 12764
rect 7156 12724 7162 12736
rect 9674 12724 9680 12776
rect 9732 12724 9738 12776
rect 9953 12767 10011 12773
rect 9953 12733 9965 12767
rect 9999 12733 10011 12767
rect 9953 12727 10011 12733
rect 3694 12656 3700 12708
rect 3752 12696 3758 12708
rect 3752 12668 6316 12696
rect 3752 12656 3758 12668
rect 3510 12588 3516 12640
rect 3568 12628 3574 12640
rect 3786 12628 3792 12640
rect 3568 12600 3792 12628
rect 3568 12588 3574 12600
rect 3786 12588 3792 12600
rect 3844 12588 3850 12640
rect 4614 12588 4620 12640
rect 4672 12588 4678 12640
rect 6288 12628 6316 12668
rect 6362 12656 6368 12708
rect 6420 12696 6426 12708
rect 6730 12696 6736 12708
rect 6420 12668 6736 12696
rect 6420 12656 6426 12668
rect 6730 12656 6736 12668
rect 6788 12656 6794 12708
rect 6932 12696 6960 12724
rect 9968 12696 9996 12727
rect 10413 12699 10471 12705
rect 10413 12696 10425 12699
rect 6932 12668 9674 12696
rect 9968 12668 10425 12696
rect 9493 12631 9551 12637
rect 9493 12628 9505 12631
rect 6288 12600 9505 12628
rect 9493 12597 9505 12600
rect 9539 12597 9551 12631
rect 9646 12628 9674 12668
rect 10413 12665 10425 12668
rect 10459 12665 10471 12699
rect 10612 12696 10640 12804
rect 10778 12792 10784 12844
rect 10836 12792 10842 12844
rect 11606 12832 11612 12844
rect 10980 12804 11612 12832
rect 10689 12767 10747 12773
rect 10689 12733 10701 12767
rect 10735 12764 10747 12767
rect 10980 12764 11008 12804
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 11793 12835 11851 12841
rect 11793 12801 11805 12835
rect 11839 12801 11851 12835
rect 11793 12795 11851 12801
rect 10735 12736 11008 12764
rect 10735 12733 10747 12736
rect 10689 12727 10747 12733
rect 11514 12724 11520 12776
rect 11572 12724 11578 12776
rect 11330 12696 11336 12708
rect 10612 12668 11336 12696
rect 10413 12659 10471 12665
rect 11330 12656 11336 12668
rect 11388 12656 11394 12708
rect 11808 12696 11836 12795
rect 11882 12792 11888 12844
rect 11940 12792 11946 12844
rect 11974 12792 11980 12844
rect 12032 12832 12038 12844
rect 12710 12832 12716 12844
rect 12032 12804 12716 12832
rect 12032 12792 12038 12804
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 13078 12792 13084 12844
rect 13136 12792 13142 12844
rect 13280 12841 13308 12872
rect 13265 12835 13323 12841
rect 13265 12801 13277 12835
rect 13311 12801 13323 12835
rect 13265 12795 13323 12801
rect 13354 12792 13360 12844
rect 13412 12832 13418 12844
rect 13633 12835 13691 12841
rect 13633 12832 13645 12835
rect 13412 12804 13645 12832
rect 13412 12792 13418 12804
rect 13633 12801 13645 12804
rect 13679 12801 13691 12835
rect 13633 12795 13691 12801
rect 12161 12767 12219 12773
rect 12161 12733 12173 12767
rect 12207 12764 12219 12767
rect 12250 12764 12256 12776
rect 12207 12736 12256 12764
rect 12207 12733 12219 12736
rect 12161 12727 12219 12733
rect 12250 12724 12256 12736
rect 12308 12724 12314 12776
rect 13096 12764 13124 12792
rect 13449 12767 13507 12773
rect 13449 12764 13461 12767
rect 13096 12736 13461 12764
rect 13449 12733 13461 12736
rect 13495 12733 13507 12767
rect 13449 12727 13507 12733
rect 13541 12767 13599 12773
rect 13541 12733 13553 12767
rect 13587 12733 13599 12767
rect 13541 12727 13599 12733
rect 11885 12699 11943 12705
rect 11885 12696 11897 12699
rect 11808 12668 11897 12696
rect 11885 12665 11897 12668
rect 11931 12665 11943 12699
rect 11885 12659 11943 12665
rect 12342 12656 12348 12708
rect 12400 12696 12406 12708
rect 13556 12696 13584 12727
rect 12400 12668 13584 12696
rect 13648 12696 13676 12795
rect 13722 12792 13728 12844
rect 13780 12792 13786 12844
rect 13832 12764 13860 12872
rect 14550 12860 14556 12912
rect 14608 12900 14614 12912
rect 14645 12903 14703 12909
rect 14645 12900 14657 12903
rect 14608 12872 14657 12900
rect 14608 12860 14614 12872
rect 14645 12869 14657 12872
rect 14691 12869 14703 12903
rect 14645 12863 14703 12869
rect 14829 12903 14887 12909
rect 14829 12869 14841 12903
rect 14875 12900 14887 12903
rect 15010 12900 15016 12912
rect 14875 12872 15016 12900
rect 14875 12869 14887 12872
rect 14829 12863 14887 12869
rect 15010 12860 15016 12872
rect 15068 12900 15074 12912
rect 15948 12900 15976 12931
rect 17310 12928 17316 12980
rect 17368 12968 17374 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 17368 12940 17785 12968
rect 17368 12928 17374 12940
rect 17773 12937 17785 12940
rect 17819 12937 17831 12971
rect 17773 12931 17831 12937
rect 15068 12872 15976 12900
rect 15068 12860 15074 12872
rect 14185 12835 14243 12841
rect 14185 12801 14197 12835
rect 14231 12832 14243 12835
rect 14274 12832 14280 12844
rect 14231 12804 14280 12832
rect 14231 12801 14243 12804
rect 14185 12795 14243 12801
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 14369 12835 14427 12841
rect 14369 12801 14381 12835
rect 14415 12832 14427 12835
rect 14458 12832 14464 12844
rect 14415 12804 14464 12832
rect 14415 12801 14427 12804
rect 14369 12795 14427 12801
rect 14458 12792 14464 12804
rect 14516 12792 14522 12844
rect 14734 12792 14740 12844
rect 14792 12832 14798 12844
rect 15304 12841 15332 12872
rect 16390 12860 16396 12912
rect 16448 12900 16454 12912
rect 16448 12872 16712 12900
rect 16448 12860 16454 12872
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 14792 12804 14933 12832
rect 14792 12792 14798 12804
rect 14921 12801 14933 12804
rect 14967 12801 14979 12835
rect 14921 12795 14979 12801
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12801 15347 12835
rect 15289 12795 15347 12801
rect 15565 12835 15623 12841
rect 15565 12801 15577 12835
rect 15611 12832 15623 12835
rect 15746 12832 15752 12844
rect 15611 12804 15752 12832
rect 15611 12801 15623 12804
rect 15565 12795 15623 12801
rect 15746 12792 15752 12804
rect 15804 12792 15810 12844
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12801 15899 12835
rect 15841 12795 15899 12801
rect 15105 12767 15163 12773
rect 15105 12764 15117 12767
rect 13832 12736 15117 12764
rect 15105 12733 15117 12736
rect 15151 12733 15163 12767
rect 15856 12764 15884 12795
rect 16114 12792 16120 12844
rect 16172 12792 16178 12844
rect 16298 12792 16304 12844
rect 16356 12832 16362 12844
rect 16684 12841 16712 12872
rect 16485 12835 16543 12841
rect 16485 12832 16497 12835
rect 16356 12804 16497 12832
rect 16356 12792 16362 12804
rect 16485 12801 16497 12804
rect 16531 12801 16543 12835
rect 16485 12795 16543 12801
rect 16669 12835 16727 12841
rect 16669 12801 16681 12835
rect 16715 12801 16727 12835
rect 16669 12795 16727 12801
rect 17218 12792 17224 12844
rect 17276 12832 17282 12844
rect 17313 12835 17371 12841
rect 17313 12832 17325 12835
rect 17276 12804 17325 12832
rect 17276 12792 17282 12804
rect 17313 12801 17325 12804
rect 17359 12832 17371 12835
rect 17589 12835 17647 12841
rect 17589 12832 17601 12835
rect 17359 12804 17601 12832
rect 17359 12801 17371 12804
rect 17313 12795 17371 12801
rect 17589 12801 17601 12804
rect 17635 12832 17647 12835
rect 17681 12835 17739 12841
rect 17681 12832 17693 12835
rect 17635 12804 17693 12832
rect 17635 12801 17647 12804
rect 17589 12795 17647 12801
rect 17681 12801 17693 12804
rect 17727 12801 17739 12835
rect 17681 12795 17739 12801
rect 16316 12764 16344 12792
rect 15856 12736 16344 12764
rect 15105 12727 15163 12733
rect 14277 12699 14335 12705
rect 14277 12696 14289 12699
rect 13648 12668 14289 12696
rect 12400 12656 12406 12668
rect 14277 12665 14289 12668
rect 14323 12665 14335 12699
rect 14277 12659 14335 12665
rect 14826 12656 14832 12708
rect 14884 12696 14890 12708
rect 15010 12696 15016 12708
rect 14884 12668 15016 12696
rect 14884 12656 14890 12668
rect 15010 12656 15016 12668
rect 15068 12656 15074 12708
rect 16390 12656 16396 12708
rect 16448 12696 16454 12708
rect 17221 12699 17279 12705
rect 17221 12696 17233 12699
rect 16448 12668 17233 12696
rect 16448 12656 16454 12668
rect 17221 12665 17233 12668
rect 17267 12665 17279 12699
rect 17221 12659 17279 12665
rect 10686 12628 10692 12640
rect 9646 12600 10692 12628
rect 9493 12591 9551 12597
rect 10686 12588 10692 12600
rect 10744 12588 10750 12640
rect 10781 12631 10839 12637
rect 10781 12597 10793 12631
rect 10827 12628 10839 12631
rect 11054 12628 11060 12640
rect 10827 12600 11060 12628
rect 10827 12597 10839 12600
rect 10781 12591 10839 12597
rect 11054 12588 11060 12600
rect 11112 12628 11118 12640
rect 11422 12628 11428 12640
rect 11112 12600 11428 12628
rect 11112 12588 11118 12600
rect 11422 12588 11428 12600
rect 11480 12588 11486 12640
rect 11701 12631 11759 12637
rect 11701 12597 11713 12631
rect 11747 12628 11759 12631
rect 13170 12628 13176 12640
rect 11747 12600 13176 12628
rect 11747 12597 11759 12600
rect 11701 12591 11759 12597
rect 13170 12588 13176 12600
rect 13228 12588 13234 12640
rect 13906 12588 13912 12640
rect 13964 12588 13970 12640
rect 13998 12588 14004 12640
rect 14056 12628 14062 12640
rect 14458 12628 14464 12640
rect 14056 12600 14464 12628
rect 14056 12588 14062 12600
rect 14458 12588 14464 12600
rect 14516 12628 14522 12640
rect 14645 12631 14703 12637
rect 14645 12628 14657 12631
rect 14516 12600 14657 12628
rect 14516 12588 14522 12600
rect 14645 12597 14657 12600
rect 14691 12597 14703 12631
rect 14645 12591 14703 12597
rect 15838 12588 15844 12640
rect 15896 12628 15902 12640
rect 16117 12631 16175 12637
rect 16117 12628 16129 12631
rect 15896 12600 16129 12628
rect 15896 12588 15902 12600
rect 16117 12597 16129 12600
rect 16163 12597 16175 12631
rect 16117 12591 16175 12597
rect 16206 12588 16212 12640
rect 16264 12628 16270 12640
rect 16853 12631 16911 12637
rect 16853 12628 16865 12631
rect 16264 12600 16865 12628
rect 16264 12588 16270 12600
rect 16853 12597 16865 12600
rect 16899 12597 16911 12631
rect 16853 12591 16911 12597
rect 17494 12588 17500 12640
rect 17552 12588 17558 12640
rect 1104 12538 18400 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 18400 12538
rect 1104 12464 18400 12486
rect 2409 12427 2467 12433
rect 2409 12393 2421 12427
rect 2455 12424 2467 12427
rect 2958 12424 2964 12436
rect 2455 12396 2964 12424
rect 2455 12393 2467 12396
rect 2409 12387 2467 12393
rect 2958 12384 2964 12396
rect 3016 12384 3022 12436
rect 3878 12384 3884 12436
rect 3936 12424 3942 12436
rect 3973 12427 4031 12433
rect 3973 12424 3985 12427
rect 3936 12396 3985 12424
rect 3936 12384 3942 12396
rect 3973 12393 3985 12396
rect 4019 12393 4031 12427
rect 3973 12387 4031 12393
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4249 12427 4307 12433
rect 4249 12424 4261 12427
rect 4212 12396 4261 12424
rect 4212 12384 4218 12396
rect 4249 12393 4261 12396
rect 4295 12393 4307 12427
rect 4249 12387 4307 12393
rect 5552 12396 5948 12424
rect 3326 12316 3332 12368
rect 3384 12356 3390 12368
rect 4062 12356 4068 12368
rect 3384 12328 4068 12356
rect 3384 12316 3390 12328
rect 4062 12316 4068 12328
rect 4120 12356 4126 12368
rect 4614 12356 4620 12368
rect 4120 12328 4620 12356
rect 4120 12316 4126 12328
rect 4614 12316 4620 12328
rect 4672 12316 4678 12368
rect 5552 12356 5580 12396
rect 5920 12368 5948 12396
rect 6730 12384 6736 12436
rect 6788 12384 6794 12436
rect 6840 12396 7328 12424
rect 5185 12328 5580 12356
rect 3878 12288 3884 12300
rect 2608 12260 3884 12288
rect 2608 12229 2636 12260
rect 3878 12248 3884 12260
rect 3936 12248 3942 12300
rect 4522 12248 4528 12300
rect 4580 12248 4586 12300
rect 2593 12223 2651 12229
rect 2593 12189 2605 12223
rect 2639 12189 2651 12223
rect 2593 12183 2651 12189
rect 2958 12180 2964 12232
rect 3016 12180 3022 12232
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12220 3111 12223
rect 3234 12220 3240 12232
rect 3099 12192 3240 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 3234 12180 3240 12192
rect 3292 12180 3298 12232
rect 4430 12180 4436 12232
rect 4488 12180 4494 12232
rect 4540 12220 4568 12248
rect 4801 12223 4859 12229
rect 4801 12220 4813 12223
rect 4540 12192 4813 12220
rect 4801 12189 4813 12192
rect 4847 12189 4859 12223
rect 4801 12183 4859 12189
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12220 4951 12223
rect 5185 12220 5213 12328
rect 5718 12316 5724 12368
rect 5776 12316 5782 12368
rect 5902 12316 5908 12368
rect 5960 12356 5966 12368
rect 6840 12356 6868 12396
rect 5960 12328 6868 12356
rect 6917 12359 6975 12365
rect 5960 12316 5966 12328
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 5813 12291 5871 12297
rect 5813 12288 5825 12291
rect 5592 12260 5825 12288
rect 5592 12248 5598 12260
rect 5813 12257 5825 12260
rect 5859 12288 5871 12291
rect 6362 12288 6368 12300
rect 5859 12260 6368 12288
rect 5859 12257 5871 12260
rect 5813 12251 5871 12257
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 6656 12297 6684 12328
rect 6917 12325 6929 12359
rect 6963 12356 6975 12359
rect 7190 12356 7196 12368
rect 6963 12328 7196 12356
rect 6963 12325 6975 12328
rect 6917 12319 6975 12325
rect 7190 12316 7196 12328
rect 7248 12316 7254 12368
rect 7300 12356 7328 12396
rect 7742 12384 7748 12436
rect 7800 12384 7806 12436
rect 7834 12384 7840 12436
rect 7892 12424 7898 12436
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 7892 12396 8585 12424
rect 7892 12384 7898 12396
rect 8573 12393 8585 12396
rect 8619 12393 8631 12427
rect 8573 12387 8631 12393
rect 9585 12427 9643 12433
rect 9585 12393 9597 12427
rect 9631 12424 9643 12427
rect 9858 12424 9864 12436
rect 9631 12396 9864 12424
rect 9631 12393 9643 12396
rect 9585 12387 9643 12393
rect 9858 12384 9864 12396
rect 9916 12424 9922 12436
rect 10318 12424 10324 12436
rect 9916 12396 10324 12424
rect 9916 12384 9922 12396
rect 10318 12384 10324 12396
rect 10376 12384 10382 12436
rect 11241 12427 11299 12433
rect 11241 12393 11253 12427
rect 11287 12424 11299 12427
rect 11333 12427 11391 12433
rect 11333 12424 11345 12427
rect 11287 12396 11345 12424
rect 11287 12393 11299 12396
rect 11241 12387 11299 12393
rect 11333 12393 11345 12396
rect 11379 12393 11391 12427
rect 11333 12387 11391 12393
rect 11514 12384 11520 12436
rect 11572 12424 11578 12436
rect 11793 12427 11851 12433
rect 11793 12424 11805 12427
rect 11572 12396 11805 12424
rect 11572 12384 11578 12396
rect 11793 12393 11805 12396
rect 11839 12393 11851 12427
rect 12897 12427 12955 12433
rect 11793 12387 11851 12393
rect 11993 12396 12296 12424
rect 7300 12328 7880 12356
rect 6641 12291 6699 12297
rect 6641 12257 6653 12291
rect 6687 12257 6699 12291
rect 6641 12251 6699 12257
rect 6730 12248 6736 12300
rect 6788 12288 6794 12300
rect 7852 12288 7880 12328
rect 8294 12316 8300 12368
rect 8352 12356 8358 12368
rect 8478 12356 8484 12368
rect 8352 12328 8484 12356
rect 8352 12316 8358 12328
rect 8478 12316 8484 12328
rect 8536 12316 8542 12368
rect 8680 12328 9352 12356
rect 8680 12288 8708 12328
rect 6788 12260 7788 12288
rect 7852 12260 8708 12288
rect 6788 12248 6794 12260
rect 4939 12192 5213 12220
rect 5261 12223 5319 12229
rect 4939 12189 4951 12192
rect 4893 12183 4951 12189
rect 5261 12189 5273 12223
rect 5307 12189 5319 12223
rect 5261 12183 5319 12189
rect 2685 12155 2743 12161
rect 2685 12121 2697 12155
rect 2731 12121 2743 12155
rect 2685 12115 2743 12121
rect 2777 12155 2835 12161
rect 2777 12121 2789 12155
rect 2823 12152 2835 12155
rect 3418 12152 3424 12164
rect 2823 12124 3424 12152
rect 2823 12121 2835 12124
rect 2777 12115 2835 12121
rect 2700 12084 2728 12115
rect 3418 12112 3424 12124
rect 3476 12152 3482 12164
rect 3789 12155 3847 12161
rect 3789 12152 3801 12155
rect 3476 12124 3801 12152
rect 3476 12112 3482 12124
rect 3789 12121 3801 12124
rect 3835 12121 3847 12155
rect 3789 12115 3847 12121
rect 3878 12112 3884 12164
rect 3936 12152 3942 12164
rect 4525 12155 4583 12161
rect 4525 12152 4537 12155
rect 3936 12124 4537 12152
rect 3936 12112 3942 12124
rect 4525 12121 4537 12124
rect 4571 12121 4583 12155
rect 4525 12115 4583 12121
rect 4614 12112 4620 12164
rect 4672 12152 4678 12164
rect 5276 12152 5304 12183
rect 5442 12180 5448 12232
rect 5500 12180 5506 12232
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12220 6607 12223
rect 7098 12220 7104 12232
rect 6595 12192 7104 12220
rect 6595 12189 6607 12192
rect 6549 12183 6607 12189
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 7190 12180 7196 12232
rect 7248 12180 7254 12232
rect 7282 12180 7288 12232
rect 7340 12180 7346 12232
rect 7374 12180 7380 12232
rect 7432 12180 7438 12232
rect 7466 12180 7472 12232
rect 7524 12180 7530 12232
rect 7653 12223 7711 12229
rect 7653 12189 7665 12223
rect 7699 12189 7711 12223
rect 7653 12183 7711 12189
rect 7668 12152 7696 12183
rect 4672 12124 5304 12152
rect 6932 12124 7696 12152
rect 7760 12152 7788 12260
rect 8754 12248 8760 12300
rect 8812 12288 8818 12300
rect 9324 12288 9352 12328
rect 9674 12316 9680 12368
rect 9732 12356 9738 12368
rect 10594 12356 10600 12368
rect 9732 12328 10600 12356
rect 9732 12316 9738 12328
rect 10594 12316 10600 12328
rect 10652 12316 10658 12368
rect 11993 12356 12021 12396
rect 10704 12328 12021 12356
rect 9950 12288 9956 12300
rect 8812 12260 9260 12288
rect 9324 12260 9956 12288
rect 8812 12248 8818 12260
rect 7834 12180 7840 12232
rect 7892 12220 7898 12232
rect 7929 12223 7987 12229
rect 7929 12220 7941 12223
rect 7892 12192 7941 12220
rect 7892 12180 7898 12192
rect 7929 12189 7941 12192
rect 7975 12189 7987 12223
rect 7929 12183 7987 12189
rect 8018 12180 8024 12232
rect 8076 12220 8082 12232
rect 8297 12223 8355 12229
rect 8297 12220 8309 12223
rect 8076 12192 8309 12220
rect 8076 12180 8082 12192
rect 8297 12189 8309 12192
rect 8343 12220 8355 12223
rect 8404 12220 8616 12222
rect 8846 12220 8852 12232
rect 8343 12194 8852 12220
rect 8343 12192 8432 12194
rect 8588 12192 8852 12194
rect 8343 12189 8355 12192
rect 8297 12183 8355 12189
rect 8846 12180 8852 12192
rect 8904 12180 8910 12232
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 9232 12220 9260 12260
rect 9950 12248 9956 12260
rect 10008 12288 10014 12300
rect 10226 12288 10232 12300
rect 10008 12260 10232 12288
rect 10008 12248 10014 12260
rect 10226 12248 10232 12260
rect 10284 12248 10290 12300
rect 9309 12223 9367 12229
rect 9309 12220 9321 12223
rect 9232 12192 9321 12220
rect 9309 12189 9321 12192
rect 9355 12220 9367 12223
rect 10502 12220 10508 12232
rect 9355 12192 10508 12220
rect 9355 12189 9367 12192
rect 9309 12183 9367 12189
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 7760 12124 8432 12152
rect 4672 12112 4678 12124
rect 2866 12084 2872 12096
rect 2700 12056 2872 12084
rect 2866 12044 2872 12056
rect 2924 12044 2930 12096
rect 3510 12044 3516 12096
rect 3568 12084 3574 12096
rect 3989 12087 4047 12093
rect 3989 12084 4001 12087
rect 3568 12056 4001 12084
rect 3568 12044 3574 12056
rect 3989 12053 4001 12056
rect 4035 12053 4047 12087
rect 3989 12047 4047 12053
rect 4157 12087 4215 12093
rect 4157 12053 4169 12087
rect 4203 12084 4215 12087
rect 5350 12084 5356 12096
rect 4203 12056 5356 12084
rect 4203 12053 4215 12056
rect 4157 12047 4215 12053
rect 5350 12044 5356 12056
rect 5408 12084 5414 12096
rect 6932 12084 6960 12124
rect 5408 12056 6960 12084
rect 7009 12087 7067 12093
rect 5408 12044 5414 12056
rect 7009 12053 7021 12087
rect 7055 12084 7067 12087
rect 7190 12084 7196 12096
rect 7055 12056 7196 12084
rect 7055 12053 7067 12056
rect 7009 12047 7067 12053
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 7742 12044 7748 12096
rect 7800 12084 7806 12096
rect 8404 12093 8432 12124
rect 8570 12112 8576 12164
rect 8628 12112 8634 12164
rect 9677 12155 9735 12161
rect 8680 12124 9536 12152
rect 8205 12087 8263 12093
rect 8205 12084 8217 12087
rect 7800 12056 8217 12084
rect 7800 12044 7806 12056
rect 8205 12053 8217 12056
rect 8251 12053 8263 12087
rect 8205 12047 8263 12053
rect 8389 12087 8447 12093
rect 8389 12053 8401 12087
rect 8435 12084 8447 12087
rect 8680 12084 8708 12124
rect 8435 12056 8708 12084
rect 8435 12053 8447 12056
rect 8389 12047 8447 12053
rect 9122 12044 9128 12096
rect 9180 12084 9186 12096
rect 9398 12084 9404 12096
rect 9180 12056 9404 12084
rect 9180 12044 9186 12056
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 9508 12084 9536 12124
rect 9677 12121 9689 12155
rect 9723 12152 9735 12155
rect 10042 12152 10048 12164
rect 9723 12124 10048 12152
rect 9723 12121 9735 12124
rect 9677 12115 9735 12121
rect 10042 12112 10048 12124
rect 10100 12112 10106 12164
rect 10704 12084 10732 12328
rect 10870 12248 10876 12300
rect 10928 12288 10934 12300
rect 10928 12260 11376 12288
rect 10928 12248 10934 12260
rect 11054 12180 11060 12232
rect 11112 12180 11118 12232
rect 11238 12180 11244 12232
rect 11296 12180 11302 12232
rect 11348 12220 11376 12260
rect 11422 12248 11428 12300
rect 11480 12248 11486 12300
rect 11609 12223 11667 12229
rect 11609 12220 11621 12223
rect 11348 12192 11621 12220
rect 11609 12189 11621 12192
rect 11655 12189 11667 12223
rect 11609 12183 11667 12189
rect 11698 12180 11704 12232
rect 11756 12220 11762 12232
rect 11885 12223 11943 12229
rect 11885 12220 11897 12223
rect 11756 12192 11897 12220
rect 11756 12180 11762 12192
rect 11885 12189 11897 12192
rect 11931 12189 11943 12223
rect 11885 12183 11943 12189
rect 12069 12223 12127 12229
rect 12069 12189 12081 12223
rect 12115 12189 12127 12223
rect 12069 12183 12127 12189
rect 10778 12112 10784 12164
rect 10836 12152 10842 12164
rect 11333 12155 11391 12161
rect 11333 12152 11345 12155
rect 10836 12124 11345 12152
rect 10836 12112 10842 12124
rect 11333 12121 11345 12124
rect 11379 12121 11391 12155
rect 11333 12115 11391 12121
rect 11422 12112 11428 12164
rect 11480 12152 11486 12164
rect 12084 12152 12112 12183
rect 11480 12124 12112 12152
rect 12268 12152 12296 12396
rect 12897 12393 12909 12427
rect 12943 12424 12955 12427
rect 13446 12424 13452 12436
rect 12943 12396 13452 12424
rect 12943 12393 12955 12396
rect 12897 12387 12955 12393
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 13556 12396 14688 12424
rect 13556 12356 13584 12396
rect 12820 12328 13584 12356
rect 12342 12180 12348 12232
rect 12400 12220 12406 12232
rect 12621 12223 12679 12229
rect 12621 12220 12633 12223
rect 12400 12192 12633 12220
rect 12400 12180 12406 12192
rect 12621 12189 12633 12192
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 12713 12223 12771 12229
rect 12713 12189 12725 12223
rect 12759 12220 12771 12223
rect 12820 12220 12848 12328
rect 13722 12316 13728 12368
rect 13780 12316 13786 12368
rect 14182 12316 14188 12368
rect 14240 12356 14246 12368
rect 14550 12356 14556 12368
rect 14240 12328 14556 12356
rect 14240 12316 14246 12328
rect 14550 12316 14556 12328
rect 14608 12316 14614 12368
rect 14660 12356 14688 12396
rect 15194 12384 15200 12436
rect 15252 12424 15258 12436
rect 15565 12427 15623 12433
rect 15565 12424 15577 12427
rect 15252 12396 15577 12424
rect 15252 12384 15258 12396
rect 15565 12393 15577 12396
rect 15611 12393 15623 12427
rect 15565 12387 15623 12393
rect 15930 12384 15936 12436
rect 15988 12384 15994 12436
rect 15654 12356 15660 12368
rect 14660 12328 15660 12356
rect 15654 12316 15660 12328
rect 15712 12316 15718 12368
rect 13449 12291 13507 12297
rect 13449 12288 13461 12291
rect 12912 12260 13461 12288
rect 12912 12229 12940 12260
rect 13449 12257 13461 12260
rect 13495 12288 13507 12291
rect 13740 12288 13768 12316
rect 16206 12288 16212 12300
rect 13495 12260 13768 12288
rect 14293 12260 16212 12288
rect 13495 12257 13507 12260
rect 13449 12251 13507 12257
rect 12759 12192 12848 12220
rect 12897 12223 12955 12229
rect 12759 12189 12771 12192
rect 12713 12183 12771 12189
rect 12897 12189 12909 12223
rect 12943 12189 12955 12223
rect 12897 12183 12955 12189
rect 13170 12180 13176 12232
rect 13228 12180 13234 12232
rect 13354 12180 13360 12232
rect 13412 12180 13418 12232
rect 13538 12180 13544 12232
rect 13596 12180 13602 12232
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 12268 12124 13216 12152
rect 11480 12112 11486 12124
rect 9508 12056 10732 12084
rect 11238 12044 11244 12096
rect 11296 12084 11302 12096
rect 11514 12084 11520 12096
rect 11296 12056 11520 12084
rect 11296 12044 11302 12056
rect 11514 12044 11520 12056
rect 11572 12044 11578 12096
rect 12069 12087 12127 12093
rect 12069 12053 12081 12087
rect 12115 12084 12127 12087
rect 12342 12084 12348 12096
rect 12115 12056 12348 12084
rect 12115 12053 12127 12056
rect 12069 12047 12127 12053
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 12986 12044 12992 12096
rect 13044 12044 13050 12096
rect 13188 12084 13216 12124
rect 13262 12112 13268 12164
rect 13320 12152 13326 12164
rect 13740 12152 13768 12183
rect 13320 12124 13768 12152
rect 13320 12112 13326 12124
rect 14293 12084 14321 12260
rect 16206 12248 16212 12260
rect 16264 12248 16270 12300
rect 14366 12180 14372 12232
rect 14424 12180 14430 12232
rect 14458 12180 14464 12232
rect 14516 12180 14522 12232
rect 14645 12223 14703 12229
rect 14645 12220 14657 12223
rect 14568 12192 14657 12220
rect 13188 12056 14321 12084
rect 14458 12044 14464 12096
rect 14516 12084 14522 12096
rect 14568 12084 14596 12192
rect 14645 12189 14657 12192
rect 14691 12189 14703 12223
rect 14645 12183 14703 12189
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12220 14795 12223
rect 14826 12220 14832 12232
rect 14783 12192 14832 12220
rect 14783 12189 14795 12192
rect 14737 12183 14795 12189
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 15105 12223 15163 12229
rect 15105 12189 15117 12223
rect 15151 12189 15163 12223
rect 15473 12223 15531 12229
rect 15473 12220 15485 12223
rect 15105 12183 15163 12189
rect 15212 12192 15485 12220
rect 15120 12152 15148 12183
rect 14660 12124 15148 12152
rect 14660 12096 14688 12124
rect 14516 12056 14596 12084
rect 14516 12044 14522 12056
rect 14642 12044 14648 12096
rect 14700 12044 14706 12096
rect 14826 12044 14832 12096
rect 14884 12084 14890 12096
rect 14921 12087 14979 12093
rect 14921 12084 14933 12087
rect 14884 12056 14933 12084
rect 14884 12044 14890 12056
rect 14921 12053 14933 12056
rect 14967 12053 14979 12087
rect 14921 12047 14979 12053
rect 15010 12044 15016 12096
rect 15068 12084 15074 12096
rect 15212 12084 15240 12192
rect 15473 12189 15485 12192
rect 15519 12189 15531 12223
rect 15473 12183 15531 12189
rect 15657 12223 15715 12229
rect 15657 12189 15669 12223
rect 15703 12189 15715 12223
rect 15657 12183 15715 12189
rect 15672 12152 15700 12183
rect 17678 12180 17684 12232
rect 17736 12180 17742 12232
rect 15304 12124 15700 12152
rect 15304 12096 15332 12124
rect 16390 12112 16396 12164
rect 16448 12112 16454 12164
rect 17310 12112 17316 12164
rect 17368 12152 17374 12164
rect 17405 12155 17463 12161
rect 17405 12152 17417 12155
rect 17368 12124 17417 12152
rect 17368 12112 17374 12124
rect 17405 12121 17417 12124
rect 17451 12121 17463 12155
rect 17405 12115 17463 12121
rect 15068 12056 15240 12084
rect 15068 12044 15074 12056
rect 15286 12044 15292 12096
rect 15344 12044 15350 12096
rect 1104 11994 18400 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 18400 11994
rect 1104 11920 18400 11942
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3053 11883 3111 11889
rect 3053 11880 3065 11883
rect 3016 11852 3065 11880
rect 3016 11840 3022 11852
rect 3053 11849 3065 11852
rect 3099 11849 3111 11883
rect 3053 11843 3111 11849
rect 3234 11840 3240 11892
rect 3292 11880 3298 11892
rect 4341 11883 4399 11889
rect 3292 11852 4108 11880
rect 3292 11840 3298 11852
rect 3510 11772 3516 11824
rect 3568 11812 3574 11824
rect 3973 11815 4031 11821
rect 3973 11812 3985 11815
rect 3568 11784 3985 11812
rect 3568 11772 3574 11784
rect 3973 11781 3985 11784
rect 4019 11781 4031 11815
rect 4080 11812 4108 11852
rect 4341 11849 4353 11883
rect 4387 11880 4399 11883
rect 4430 11880 4436 11892
rect 4387 11852 4436 11880
rect 4387 11849 4399 11852
rect 4341 11843 4399 11849
rect 4430 11840 4436 11852
rect 4488 11880 4494 11892
rect 6454 11880 6460 11892
rect 4488 11852 6460 11880
rect 4488 11840 4494 11852
rect 6454 11840 6460 11852
rect 6512 11840 6518 11892
rect 7190 11840 7196 11892
rect 7248 11840 7254 11892
rect 7374 11840 7380 11892
rect 7432 11880 7438 11892
rect 7837 11883 7895 11889
rect 7837 11880 7849 11883
rect 7432 11852 7849 11880
rect 7432 11840 7438 11852
rect 7837 11849 7849 11852
rect 7883 11849 7895 11883
rect 7837 11843 7895 11849
rect 8496 11852 10364 11880
rect 5534 11812 5540 11824
rect 4080 11784 5540 11812
rect 3973 11775 4031 11781
rect 5534 11772 5540 11784
rect 5592 11772 5598 11824
rect 5902 11772 5908 11824
rect 5960 11812 5966 11824
rect 7558 11812 7564 11824
rect 5960 11784 7564 11812
rect 5960 11772 5966 11784
rect 7558 11772 7564 11784
rect 7616 11772 7622 11824
rect 7653 11815 7711 11821
rect 7653 11781 7665 11815
rect 7699 11812 7711 11815
rect 8496 11812 8524 11852
rect 7699 11784 8524 11812
rect 7699 11781 7711 11784
rect 7653 11775 7711 11781
rect 8938 11772 8944 11824
rect 8996 11812 9002 11824
rect 9585 11815 9643 11821
rect 9585 11812 9597 11815
rect 8996 11784 9597 11812
rect 8996 11772 9002 11784
rect 9585 11781 9597 11784
rect 9631 11781 9643 11815
rect 9585 11775 9643 11781
rect 9677 11815 9735 11821
rect 9677 11781 9689 11815
rect 9723 11781 9735 11815
rect 10336 11812 10364 11852
rect 10502 11840 10508 11892
rect 10560 11880 10566 11892
rect 12989 11883 13047 11889
rect 10560 11852 12434 11880
rect 10560 11840 10566 11852
rect 11790 11812 11796 11824
rect 10336 11784 11796 11812
rect 9677 11775 9735 11781
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 2590 11744 2596 11756
rect 2455 11716 2596 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 2590 11704 2596 11716
rect 2648 11704 2654 11756
rect 2958 11704 2964 11756
rect 3016 11704 3022 11756
rect 3145 11747 3203 11753
rect 3145 11713 3157 11747
rect 3191 11744 3203 11747
rect 3418 11744 3424 11756
rect 3191 11716 3424 11744
rect 3191 11713 3203 11716
rect 3145 11707 3203 11713
rect 3418 11704 3424 11716
rect 3476 11744 3482 11756
rect 3697 11747 3755 11753
rect 3697 11744 3709 11747
rect 3476 11716 3709 11744
rect 3476 11704 3482 11716
rect 3697 11713 3709 11716
rect 3743 11713 3755 11747
rect 3697 11707 3755 11713
rect 3786 11704 3792 11756
rect 3844 11744 3850 11756
rect 3844 11716 3889 11744
rect 3844 11704 3850 11716
rect 4062 11704 4068 11756
rect 4120 11704 4126 11756
rect 4203 11747 4261 11753
rect 4203 11713 4215 11747
rect 4249 11744 4261 11747
rect 4614 11744 4620 11756
rect 4249 11716 4620 11744
rect 4249 11713 4261 11716
rect 4203 11707 4261 11713
rect 2682 11636 2688 11688
rect 2740 11636 2746 11688
rect 2777 11679 2835 11685
rect 2777 11645 2789 11679
rect 2823 11676 2835 11679
rect 2866 11676 2872 11688
rect 2823 11648 2872 11676
rect 2823 11645 2835 11648
rect 2777 11639 2835 11645
rect 2866 11636 2872 11648
rect 2924 11676 2930 11688
rect 4218 11676 4246 11707
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 8018 11704 8024 11756
rect 8076 11704 8082 11756
rect 8110 11704 8116 11756
rect 8168 11704 8174 11756
rect 8294 11704 8300 11756
rect 8352 11704 8358 11756
rect 8389 11747 8447 11753
rect 8389 11713 8401 11747
rect 8435 11744 8447 11747
rect 8662 11744 8668 11756
rect 8435 11716 8668 11744
rect 8435 11713 8447 11716
rect 8389 11707 8447 11713
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 9306 11753 9312 11756
rect 9297 11747 9312 11753
rect 9297 11713 9309 11747
rect 9297 11707 9312 11713
rect 9306 11704 9312 11707
rect 9364 11704 9370 11756
rect 9398 11704 9404 11756
rect 9456 11744 9462 11756
rect 9692 11744 9720 11775
rect 11790 11772 11796 11784
rect 11848 11772 11854 11824
rect 12406 11812 12434 11852
rect 12989 11849 13001 11883
rect 13035 11880 13047 11883
rect 13538 11880 13544 11892
rect 13035 11852 13544 11880
rect 13035 11849 13047 11852
rect 12989 11843 13047 11849
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 14642 11840 14648 11892
rect 14700 11840 14706 11892
rect 13722 11812 13728 11824
rect 12406 11784 13728 11812
rect 9456 11716 9501 11744
rect 9600 11716 9720 11744
rect 9769 11747 9827 11753
rect 9456 11704 9462 11716
rect 2924 11648 4246 11676
rect 2924 11636 2930 11648
rect 5994 11636 6000 11688
rect 6052 11676 6058 11688
rect 6730 11676 6736 11688
rect 6052 11648 6736 11676
rect 6052 11636 6058 11648
rect 6730 11636 6736 11648
rect 6788 11636 6794 11688
rect 7101 11679 7159 11685
rect 7101 11645 7113 11679
rect 7147 11676 7159 11679
rect 7558 11676 7564 11688
rect 7147 11648 7564 11676
rect 7147 11645 7159 11648
rect 7101 11639 7159 11645
rect 7558 11636 7564 11648
rect 7616 11636 7622 11688
rect 9490 11636 9496 11688
rect 9548 11676 9554 11688
rect 9600 11676 9628 11716
rect 9769 11713 9781 11747
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 10135 11750 10193 11753
rect 10318 11750 10324 11756
rect 10135 11747 10324 11750
rect 10135 11713 10147 11747
rect 10181 11722 10324 11747
rect 10181 11713 10193 11722
rect 10135 11707 10193 11713
rect 9548 11648 9628 11676
rect 9548 11636 9554 11648
rect 9674 11636 9680 11688
rect 9732 11676 9738 11688
rect 9784 11676 9812 11707
rect 9732 11648 9812 11676
rect 9732 11636 9738 11648
rect 6638 11568 6644 11620
rect 6696 11608 6702 11620
rect 7653 11611 7711 11617
rect 6696 11580 7604 11608
rect 6696 11568 6702 11580
rect 4890 11500 4896 11552
rect 4948 11540 4954 11552
rect 6730 11540 6736 11552
rect 4948 11512 6736 11540
rect 4948 11500 4954 11512
rect 6730 11500 6736 11512
rect 6788 11500 6794 11552
rect 6914 11500 6920 11552
rect 6972 11500 6978 11552
rect 7576 11540 7604 11580
rect 7653 11577 7665 11611
rect 7699 11608 7711 11611
rect 7926 11608 7932 11620
rect 7699 11580 7932 11608
rect 7699 11577 7711 11580
rect 7653 11571 7711 11577
rect 7926 11568 7932 11580
rect 7984 11568 7990 11620
rect 8110 11568 8116 11620
rect 8168 11608 8174 11620
rect 8294 11608 8300 11620
rect 8168 11580 8300 11608
rect 8168 11568 8174 11580
rect 8294 11568 8300 11580
rect 8352 11608 8358 11620
rect 8478 11608 8484 11620
rect 8352 11580 8484 11608
rect 8352 11568 8358 11580
rect 8478 11568 8484 11580
rect 8536 11568 8542 11620
rect 9309 11611 9367 11617
rect 9309 11577 9321 11611
rect 9355 11608 9367 11611
rect 9355 11580 9536 11608
rect 9355 11577 9367 11580
rect 9309 11571 9367 11577
rect 9122 11540 9128 11552
rect 7576 11512 9128 11540
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 9508 11540 9536 11580
rect 9582 11568 9588 11620
rect 9640 11608 9646 11620
rect 9766 11608 9772 11620
rect 9640 11580 9772 11608
rect 9640 11568 9646 11580
rect 9766 11568 9772 11580
rect 9824 11568 9830 11620
rect 9674 11540 9680 11552
rect 9508 11512 9680 11540
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 9858 11500 9864 11552
rect 9916 11540 9922 11552
rect 9968 11540 9996 11707
rect 10318 11704 10324 11722
rect 10376 11704 10382 11756
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 12452 11753 12480 11784
rect 13722 11772 13728 11784
rect 13780 11772 13786 11824
rect 14660 11812 14688 11840
rect 14292 11784 14688 11812
rect 12253 11747 12311 11753
rect 12253 11744 12265 11747
rect 12124 11716 12265 11744
rect 12124 11704 12130 11716
rect 12253 11713 12265 11716
rect 12299 11713 12311 11747
rect 12253 11707 12311 11713
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11713 12495 11747
rect 12437 11707 12495 11713
rect 12894 11704 12900 11756
rect 12952 11704 12958 11756
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11713 13139 11747
rect 13081 11707 13139 11713
rect 12342 11676 12348 11688
rect 10336 11648 12348 11676
rect 10336 11608 10364 11648
rect 12342 11636 12348 11648
rect 12400 11636 12406 11688
rect 13096 11676 13124 11707
rect 14090 11704 14096 11756
rect 14148 11704 14154 11756
rect 14292 11753 14320 11784
rect 14277 11747 14335 11753
rect 14277 11713 14289 11747
rect 14323 11713 14335 11747
rect 14277 11707 14335 11713
rect 14458 11704 14464 11756
rect 14516 11744 14522 11756
rect 14642 11744 14648 11756
rect 14516 11716 14648 11744
rect 14516 11704 14522 11716
rect 14642 11704 14648 11716
rect 14700 11744 14706 11756
rect 14829 11747 14887 11753
rect 14829 11744 14841 11747
rect 14700 11716 14841 11744
rect 14700 11704 14706 11716
rect 14829 11713 14841 11716
rect 14875 11713 14887 11747
rect 14829 11707 14887 11713
rect 15013 11747 15071 11753
rect 15013 11713 15025 11747
rect 15059 11713 15071 11747
rect 15013 11707 15071 11713
rect 13170 11676 13176 11688
rect 13096 11648 13176 11676
rect 13170 11636 13176 11648
rect 13228 11676 13234 11688
rect 15028 11676 15056 11707
rect 16758 11704 16764 11756
rect 16816 11744 16822 11756
rect 17954 11744 17960 11756
rect 16816 11716 17960 11744
rect 16816 11704 16822 11716
rect 17954 11704 17960 11716
rect 18012 11704 18018 11756
rect 13228 11648 15056 11676
rect 13228 11636 13234 11648
rect 10244 11580 10364 11608
rect 10244 11540 10272 11580
rect 11514 11568 11520 11620
rect 11572 11608 11578 11620
rect 12158 11608 12164 11620
rect 11572 11580 12164 11608
rect 11572 11568 11578 11580
rect 12158 11568 12164 11580
rect 12216 11568 12222 11620
rect 12526 11568 12532 11620
rect 12584 11608 12590 11620
rect 14366 11608 14372 11620
rect 12584 11580 14372 11608
rect 12584 11568 12590 11580
rect 14366 11568 14372 11580
rect 14424 11568 14430 11620
rect 14550 11568 14556 11620
rect 14608 11608 14614 11620
rect 15838 11608 15844 11620
rect 14608 11580 15844 11608
rect 14608 11568 14614 11580
rect 15838 11568 15844 11580
rect 15896 11608 15902 11620
rect 16942 11608 16948 11620
rect 15896 11580 16948 11608
rect 15896 11568 15902 11580
rect 16942 11568 16948 11580
rect 17000 11608 17006 11620
rect 17586 11608 17592 11620
rect 17000 11580 17592 11608
rect 17000 11568 17006 11580
rect 17586 11568 17592 11580
rect 17644 11568 17650 11620
rect 9916 11512 10272 11540
rect 10321 11543 10379 11549
rect 9916 11500 9922 11512
rect 10321 11509 10333 11543
rect 10367 11540 10379 11543
rect 10410 11540 10416 11552
rect 10367 11512 10416 11540
rect 10367 11509 10379 11512
rect 10321 11503 10379 11509
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 10686 11500 10692 11552
rect 10744 11540 10750 11552
rect 12250 11540 12256 11552
rect 10744 11512 12256 11540
rect 10744 11500 10750 11512
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 12710 11500 12716 11552
rect 12768 11540 12774 11552
rect 13078 11540 13084 11552
rect 12768 11512 13084 11540
rect 12768 11500 12774 11512
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 14185 11543 14243 11549
rect 14185 11540 14197 11543
rect 13872 11512 14197 11540
rect 13872 11500 13878 11512
rect 14185 11509 14197 11512
rect 14231 11509 14243 11543
rect 14185 11503 14243 11509
rect 15010 11500 15016 11552
rect 15068 11540 15074 11552
rect 15105 11543 15163 11549
rect 15105 11540 15117 11543
rect 15068 11512 15117 11540
rect 15068 11500 15074 11512
rect 15105 11509 15117 11512
rect 15151 11509 15163 11543
rect 15105 11503 15163 11509
rect 15654 11500 15660 11552
rect 15712 11540 15718 11552
rect 15930 11540 15936 11552
rect 15712 11512 15936 11540
rect 15712 11500 15718 11512
rect 15930 11500 15936 11512
rect 15988 11500 15994 11552
rect 1104 11450 18400 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 18400 11450
rect 1104 11376 18400 11398
rect 3789 11339 3847 11345
rect 3789 11305 3801 11339
rect 3835 11336 3847 11339
rect 3970 11336 3976 11348
rect 3835 11308 3976 11336
rect 3835 11305 3847 11308
rect 3789 11299 3847 11305
rect 3970 11296 3976 11308
rect 4028 11296 4034 11348
rect 4706 11296 4712 11348
rect 4764 11336 4770 11348
rect 5261 11339 5319 11345
rect 5261 11336 5273 11339
rect 4764 11308 5273 11336
rect 4764 11296 4770 11308
rect 5261 11305 5273 11308
rect 5307 11305 5319 11339
rect 6457 11339 6515 11345
rect 6457 11336 6469 11339
rect 5261 11299 5319 11305
rect 5460 11308 6469 11336
rect 4062 11268 4068 11280
rect 2516 11240 4068 11268
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11101 2007 11135
rect 1949 11095 2007 11101
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11132 2191 11135
rect 2225 11135 2283 11141
rect 2225 11132 2237 11135
rect 2179 11104 2237 11132
rect 2179 11101 2191 11104
rect 2133 11095 2191 11101
rect 2225 11101 2237 11104
rect 2271 11132 2283 11135
rect 2516 11132 2544 11240
rect 4062 11228 4068 11240
rect 4120 11228 4126 11280
rect 4157 11271 4215 11277
rect 4157 11237 4169 11271
rect 4203 11268 4215 11271
rect 4246 11268 4252 11280
rect 4203 11240 4252 11268
rect 4203 11237 4215 11240
rect 4157 11231 4215 11237
rect 4246 11228 4252 11240
rect 4304 11228 4310 11280
rect 3988 11172 5212 11200
rect 2271 11104 2544 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 1964 11064 1992 11095
rect 2590 11092 2596 11144
rect 2648 11092 2654 11144
rect 2682 11092 2688 11144
rect 2740 11132 2746 11144
rect 2869 11135 2927 11141
rect 2869 11132 2881 11135
rect 2740 11104 2881 11132
rect 2740 11092 2746 11104
rect 2869 11101 2881 11104
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 3418 11092 3424 11144
rect 3476 11132 3482 11144
rect 3988 11141 4016 11172
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3476 11104 3985 11132
rect 3476 11092 3482 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 4249 11135 4307 11141
rect 4249 11101 4261 11135
rect 4295 11101 4307 11135
rect 4249 11095 4307 11101
rect 2608 11064 2636 11092
rect 1964 11036 2636 11064
rect 2958 11024 2964 11076
rect 3016 11064 3022 11076
rect 3510 11064 3516 11076
rect 3016 11036 3516 11064
rect 3016 11024 3022 11036
rect 3510 11024 3516 11036
rect 3568 11064 3574 11076
rect 4264 11064 4292 11095
rect 4614 11092 4620 11144
rect 4672 11132 4678 11144
rect 4798 11132 4804 11144
rect 4672 11104 4804 11132
rect 4672 11092 4678 11104
rect 4798 11092 4804 11104
rect 4856 11132 4862 11144
rect 5184 11141 5212 11172
rect 5460 11141 5488 11308
rect 6457 11305 6469 11308
rect 6503 11305 6515 11339
rect 6457 11299 6515 11305
rect 7558 11296 7564 11348
rect 7616 11296 7622 11348
rect 8389 11339 8447 11345
rect 8389 11336 8401 11339
rect 7668 11308 8401 11336
rect 5718 11228 5724 11280
rect 5776 11228 5782 11280
rect 6270 11228 6276 11280
rect 6328 11228 6334 11280
rect 6730 11228 6736 11280
rect 6788 11268 6794 11280
rect 7668 11268 7696 11308
rect 8389 11305 8401 11308
rect 8435 11305 8447 11339
rect 8389 11299 8447 11305
rect 9490 11296 9496 11348
rect 9548 11336 9554 11348
rect 9548 11308 9812 11336
rect 9548 11296 9554 11308
rect 8205 11271 8263 11277
rect 8205 11268 8217 11271
rect 6788 11240 7696 11268
rect 7852 11240 8217 11268
rect 6788 11228 6794 11240
rect 4985 11135 5043 11141
rect 4985 11132 4997 11135
rect 4856 11104 4997 11132
rect 4856 11092 4862 11104
rect 4985 11101 4997 11104
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11101 5227 11135
rect 5169 11095 5227 11101
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11101 5503 11135
rect 5445 11095 5503 11101
rect 5629 11135 5687 11141
rect 5629 11101 5641 11135
rect 5675 11132 5687 11135
rect 5736 11132 5764 11228
rect 7098 11200 7104 11212
rect 6288 11172 7104 11200
rect 5675 11104 5764 11132
rect 5675 11101 5687 11104
rect 5629 11095 5687 11101
rect 5902 11092 5908 11144
rect 5960 11092 5966 11144
rect 5994 11092 6000 11144
rect 6052 11092 6058 11144
rect 6288 11141 6316 11172
rect 7098 11160 7104 11172
rect 7156 11200 7162 11212
rect 7374 11200 7380 11212
rect 7156 11172 7380 11200
rect 7156 11160 7162 11172
rect 7374 11160 7380 11172
rect 7432 11160 7438 11212
rect 7742 11160 7748 11212
rect 7800 11160 7806 11212
rect 7852 11209 7880 11240
rect 8205 11237 8217 11240
rect 8251 11237 8263 11271
rect 8205 11231 8263 11237
rect 8938 11228 8944 11280
rect 8996 11228 9002 11280
rect 7837 11203 7895 11209
rect 7837 11169 7849 11203
rect 7883 11169 7895 11203
rect 7837 11163 7895 11169
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11200 8539 11203
rect 9398 11200 9404 11212
rect 8527 11172 9404 11200
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 9398 11160 9404 11172
rect 9456 11200 9462 11212
rect 9784 11200 9812 11308
rect 10410 11296 10416 11348
rect 10468 11296 10474 11348
rect 11422 11336 11428 11348
rect 11165 11308 11428 11336
rect 9950 11228 9956 11280
rect 10008 11268 10014 11280
rect 10229 11271 10287 11277
rect 10229 11268 10241 11271
rect 10008 11240 10241 11268
rect 10008 11228 10014 11240
rect 10229 11237 10241 11240
rect 10275 11237 10287 11271
rect 10229 11231 10287 11237
rect 10686 11200 10692 11212
rect 9456 11172 9536 11200
rect 9784 11172 10692 11200
rect 9456 11160 9462 11172
rect 6273 11135 6331 11141
rect 6273 11101 6285 11135
rect 6319 11101 6331 11135
rect 6273 11095 6331 11101
rect 6638 11092 6644 11144
rect 6696 11092 6702 11144
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11132 6791 11135
rect 6822 11132 6828 11144
rect 6779 11104 6828 11132
rect 6779 11101 6791 11104
rect 6733 11095 6791 11101
rect 6822 11092 6828 11104
rect 6880 11092 6886 11144
rect 6914 11092 6920 11144
rect 6972 11092 6978 11144
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11101 7067 11135
rect 7009 11095 7067 11101
rect 4890 11064 4896 11076
rect 3568 11036 4896 11064
rect 3568 11024 3574 11036
rect 4890 11024 4896 11036
rect 4948 11024 4954 11076
rect 5074 11024 5080 11076
rect 5132 11024 5138 11076
rect 5534 11024 5540 11076
rect 5592 11024 5598 11076
rect 5810 11073 5816 11076
rect 5767 11067 5816 11073
rect 5767 11033 5779 11067
rect 5813 11033 5816 11067
rect 5767 11027 5816 11033
rect 5810 11024 5816 11027
rect 5868 11024 5874 11076
rect 6086 11024 6092 11076
rect 6144 11064 6150 11076
rect 6546 11064 6552 11076
rect 6144 11036 6552 11064
rect 6144 11024 6150 11036
rect 6546 11024 6552 11036
rect 6604 11024 6610 11076
rect 7024 11064 7052 11095
rect 7926 11092 7932 11144
rect 7984 11092 7990 11144
rect 8018 11092 8024 11144
rect 8076 11132 8082 11144
rect 8202 11132 8208 11144
rect 8076 11104 8208 11132
rect 8076 11092 8082 11104
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 8570 11092 8576 11144
rect 8628 11092 8634 11144
rect 8662 11092 8668 11144
rect 8720 11132 8726 11144
rect 9217 11135 9275 11141
rect 9217 11134 9229 11135
rect 9048 11132 9229 11134
rect 8720 11106 9229 11132
rect 8720 11104 9076 11106
rect 8720 11092 8726 11104
rect 9217 11101 9229 11106
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 7742 11064 7748 11076
rect 7024 11036 7748 11064
rect 2130 10956 2136 11008
rect 2188 10956 2194 11008
rect 3694 10956 3700 11008
rect 3752 10996 3758 11008
rect 4246 10996 4252 11008
rect 3752 10968 4252 10996
rect 3752 10956 3758 10968
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 6454 10956 6460 11008
rect 6512 10996 6518 11008
rect 7024 10996 7052 11036
rect 7742 11024 7748 11036
rect 7800 11024 7806 11076
rect 8754 11024 8760 11076
rect 8812 11064 8818 11076
rect 8941 11067 8999 11073
rect 8941 11064 8953 11067
rect 8812 11036 8953 11064
rect 8812 11024 8818 11036
rect 8941 11033 8953 11036
rect 8987 11033 8999 11067
rect 8941 11027 8999 11033
rect 9122 11024 9128 11076
rect 9180 11024 9186 11076
rect 9232 11064 9260 11095
rect 9398 11064 9404 11076
rect 9232 11036 9404 11064
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 9508 11064 9536 11172
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 9677 11135 9735 11141
rect 9677 11132 9689 11135
rect 9640 11104 9689 11132
rect 9640 11092 9646 11104
rect 9677 11101 9689 11104
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 9766 11092 9772 11144
rect 9824 11132 9830 11144
rect 10060 11141 10088 11172
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 11165 11144 11193 11308
rect 11422 11296 11428 11308
rect 11480 11296 11486 11348
rect 11790 11296 11796 11348
rect 11848 11296 11854 11348
rect 11882 11296 11888 11348
rect 11940 11336 11946 11348
rect 11940 11308 12296 11336
rect 11940 11296 11946 11308
rect 11514 11228 11520 11280
rect 11572 11228 11578 11280
rect 11701 11271 11759 11277
rect 11701 11237 11713 11271
rect 11747 11237 11759 11271
rect 11701 11231 11759 11237
rect 9861 11135 9919 11141
rect 9861 11132 9873 11135
rect 9824 11104 9873 11132
rect 9824 11092 9830 11104
rect 9861 11101 9873 11104
rect 9907 11101 9919 11135
rect 9861 11095 9919 11101
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11101 10103 11135
rect 10045 11095 10103 11101
rect 10134 11092 10140 11144
rect 10192 11092 10198 11144
rect 10870 11092 10876 11144
rect 10928 11132 10934 11144
rect 11057 11135 11115 11141
rect 11057 11132 11069 11135
rect 10928 11104 11069 11132
rect 10928 11092 10934 11104
rect 11057 11101 11069 11104
rect 11103 11101 11115 11135
rect 11057 11095 11115 11101
rect 11146 11092 11152 11144
rect 11204 11132 11210 11144
rect 11204 11104 11249 11132
rect 11204 11092 11210 11104
rect 11422 11092 11428 11144
rect 11480 11092 11486 11144
rect 11537 11141 11565 11228
rect 11716 11200 11744 11231
rect 12268 11209 12296 11308
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 14550 11336 14556 11348
rect 13044 11308 14556 11336
rect 13044 11296 13050 11308
rect 12069 11203 12127 11209
rect 12069 11200 12081 11203
rect 11716 11172 12081 11200
rect 12069 11169 12081 11172
rect 12115 11169 12127 11203
rect 12069 11163 12127 11169
rect 12253 11203 12311 11209
rect 12253 11169 12265 11203
rect 12299 11169 12311 11203
rect 12253 11163 12311 11169
rect 12342 11160 12348 11212
rect 12400 11200 12406 11212
rect 14384 11200 14412 11308
rect 14550 11296 14556 11308
rect 14608 11296 14614 11348
rect 15194 11296 15200 11348
rect 15252 11296 15258 11348
rect 17954 11296 17960 11348
rect 18012 11296 18018 11348
rect 14458 11228 14464 11280
rect 14516 11268 14522 11280
rect 14516 11240 14687 11268
rect 14516 11228 14522 11240
rect 14550 11200 14556 11212
rect 12400 11172 14320 11200
rect 14384 11172 14413 11200
rect 12400 11160 12406 11172
rect 11522 11135 11580 11141
rect 11522 11101 11534 11135
rect 11568 11101 11580 11135
rect 11522 11095 11580 11101
rect 11974 11092 11980 11144
rect 12032 11092 12038 11144
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11132 12219 11135
rect 12434 11132 12440 11144
rect 12207 11104 12440 11132
rect 12207 11101 12219 11104
rect 12161 11095 12219 11101
rect 12434 11092 12440 11104
rect 12492 11092 12498 11144
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 13633 11135 13691 11141
rect 13633 11132 13645 11135
rect 12860 11104 13645 11132
rect 12860 11092 12866 11104
rect 13633 11101 13645 11104
rect 13679 11101 13691 11135
rect 13633 11095 13691 11101
rect 13814 11092 13820 11144
rect 13872 11092 13878 11144
rect 13906 11092 13912 11144
rect 13964 11092 13970 11144
rect 14090 11092 14096 11144
rect 14148 11092 14154 11144
rect 14292 11141 14320 11172
rect 14385 11141 14413 11172
rect 14476 11172 14556 11200
rect 14476 11141 14504 11172
rect 14550 11160 14556 11172
rect 14608 11160 14614 11212
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11101 14335 11135
rect 14277 11095 14335 11101
rect 14369 11135 14427 11141
rect 14369 11101 14381 11135
rect 14415 11101 14427 11135
rect 14369 11095 14427 11101
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11101 14519 11135
rect 14659 11132 14687 11240
rect 14734 11228 14740 11280
rect 14792 11268 14798 11280
rect 14792 11240 15884 11268
rect 14792 11228 14798 11240
rect 15470 11200 15476 11212
rect 14844 11172 15476 11200
rect 14737 11135 14795 11141
rect 14737 11132 14749 11135
rect 14659 11104 14749 11132
rect 14461 11095 14519 11101
rect 14737 11101 14749 11104
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 10597 11067 10655 11073
rect 10597 11064 10609 11067
rect 9508 11036 10609 11064
rect 10597 11033 10609 11036
rect 10643 11033 10655 11067
rect 10597 11027 10655 11033
rect 11333 11067 11391 11073
rect 11333 11033 11345 11067
rect 11379 11064 11391 11067
rect 13449 11067 13507 11073
rect 11379 11036 13400 11064
rect 11379 11033 11391 11036
rect 11333 11027 11391 11033
rect 6512 10968 7052 10996
rect 6512 10956 6518 10968
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 10397 10999 10455 11005
rect 10397 10996 10409 10999
rect 8352 10968 10409 10996
rect 8352 10956 8358 10968
rect 10397 10965 10409 10968
rect 10443 10996 10455 10999
rect 10502 10996 10508 11008
rect 10443 10968 10508 10996
rect 10443 10965 10455 10968
rect 10397 10959 10455 10965
rect 10502 10956 10508 10968
rect 10560 10956 10566 11008
rect 10962 10956 10968 11008
rect 11020 10996 11026 11008
rect 12618 10996 12624 11008
rect 11020 10968 12624 10996
rect 11020 10956 11026 10968
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 13372 10996 13400 11036
rect 13449 11033 13461 11067
rect 13495 11064 13507 11067
rect 13538 11064 13544 11076
rect 13495 11036 13544 11064
rect 13495 11033 13507 11036
rect 13449 11027 13507 11033
rect 13538 11024 13544 11036
rect 13596 11024 13602 11076
rect 14599 11067 14657 11073
rect 14599 11033 14611 11067
rect 14645 11064 14657 11067
rect 14844 11064 14872 11172
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 15565 11203 15623 11209
rect 15565 11169 15577 11203
rect 15611 11200 15623 11203
rect 15746 11200 15752 11212
rect 15611 11172 15752 11200
rect 15611 11169 15623 11172
rect 15565 11163 15623 11169
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 15010 11092 15016 11144
rect 15068 11092 15074 11144
rect 15289 11135 15347 11141
rect 15289 11101 15301 11135
rect 15335 11132 15347 11135
rect 15335 11104 15608 11132
rect 15335 11101 15347 11104
rect 15289 11095 15347 11101
rect 15580 11076 15608 11104
rect 15654 11092 15660 11144
rect 15712 11092 15718 11144
rect 15856 11141 15884 11240
rect 16209 11203 16267 11209
rect 16209 11169 16221 11203
rect 16255 11200 16267 11203
rect 17678 11200 17684 11212
rect 16255 11172 17684 11200
rect 16255 11169 16267 11172
rect 16209 11163 16267 11169
rect 17678 11160 17684 11172
rect 17736 11160 17742 11212
rect 15841 11135 15899 11141
rect 15841 11101 15853 11135
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 15381 11067 15439 11073
rect 15381 11064 15393 11067
rect 14645 11036 15056 11064
rect 14645 11033 14657 11036
rect 14599 11027 14657 11033
rect 15028 11008 15056 11036
rect 15212 11036 15393 11064
rect 15212 11008 15240 11036
rect 15381 11033 15393 11036
rect 15427 11033 15439 11067
rect 15381 11027 15439 11033
rect 15562 11024 15568 11076
rect 15620 11024 15626 11076
rect 15749 11067 15807 11073
rect 15749 11033 15761 11067
rect 15795 11033 15807 11067
rect 15749 11027 15807 11033
rect 13630 10996 13636 11008
rect 13372 10968 13636 10996
rect 13630 10956 13636 10968
rect 13688 10956 13694 11008
rect 14274 10956 14280 11008
rect 14332 10996 14338 11008
rect 14829 10999 14887 11005
rect 14829 10996 14841 10999
rect 14332 10968 14841 10996
rect 14332 10956 14338 10968
rect 14829 10965 14841 10968
rect 14875 10965 14887 10999
rect 14829 10959 14887 10965
rect 15010 10956 15016 11008
rect 15068 10956 15074 11008
rect 15194 10956 15200 11008
rect 15252 10956 15258 11008
rect 15470 10956 15476 11008
rect 15528 10956 15534 11008
rect 15764 10996 15792 11027
rect 16206 11024 16212 11076
rect 16264 11064 16270 11076
rect 16485 11067 16543 11073
rect 16485 11064 16497 11067
rect 16264 11036 16497 11064
rect 16264 11024 16270 11036
rect 16485 11033 16497 11036
rect 16531 11033 16543 11067
rect 16485 11027 16543 11033
rect 17494 11024 17500 11076
rect 17552 11024 17558 11076
rect 16025 10999 16083 11005
rect 16025 10996 16037 10999
rect 15764 10968 16037 10996
rect 16025 10965 16037 10968
rect 16071 10996 16083 10999
rect 16114 10996 16120 11008
rect 16071 10968 16120 10996
rect 16071 10965 16083 10968
rect 16025 10959 16083 10965
rect 16114 10956 16120 10968
rect 16172 10956 16178 11008
rect 1104 10906 18400 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 18400 10906
rect 1104 10832 18400 10854
rect 2593 10795 2651 10801
rect 2593 10761 2605 10795
rect 2639 10792 2651 10795
rect 5442 10792 5448 10804
rect 2639 10764 4844 10792
rect 2639 10761 2651 10764
rect 2593 10755 2651 10761
rect 2866 10684 2872 10736
rect 2924 10684 2930 10736
rect 2961 10727 3019 10733
rect 2961 10693 2973 10727
rect 3007 10724 3019 10727
rect 3418 10724 3424 10736
rect 3007 10696 3424 10724
rect 3007 10693 3019 10696
rect 2961 10687 3019 10693
rect 3418 10684 3424 10696
rect 3476 10684 3482 10736
rect 3970 10684 3976 10736
rect 4028 10684 4034 10736
rect 4062 10684 4068 10736
rect 4120 10724 4126 10736
rect 4706 10724 4712 10736
rect 4120 10696 4712 10724
rect 4120 10684 4126 10696
rect 4706 10684 4712 10696
rect 4764 10684 4770 10736
rect 2130 10616 2136 10668
rect 2188 10656 2194 10668
rect 2777 10659 2835 10665
rect 2777 10656 2789 10659
rect 2188 10628 2789 10656
rect 2188 10616 2194 10628
rect 2777 10625 2789 10628
rect 2823 10625 2835 10659
rect 2777 10619 2835 10625
rect 2792 10588 2820 10619
rect 3142 10616 3148 10668
rect 3200 10616 3206 10668
rect 3234 10616 3240 10668
rect 3292 10616 3298 10668
rect 3881 10659 3939 10665
rect 3881 10625 3893 10659
rect 3927 10656 3939 10659
rect 3988 10656 4016 10684
rect 3927 10628 4016 10656
rect 3927 10625 3939 10628
rect 3881 10619 3939 10625
rect 4522 10616 4528 10668
rect 4580 10616 4586 10668
rect 4816 10665 4844 10764
rect 5184 10764 5448 10792
rect 5184 10724 5212 10764
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 5721 10795 5779 10801
rect 5721 10792 5733 10795
rect 5592 10764 5733 10792
rect 5592 10752 5598 10764
rect 5721 10761 5733 10764
rect 5767 10761 5779 10795
rect 5721 10755 5779 10761
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7009 10795 7067 10801
rect 7009 10792 7021 10795
rect 6972 10764 7021 10792
rect 6972 10752 6978 10764
rect 7009 10761 7021 10764
rect 7055 10761 7067 10795
rect 7009 10755 7067 10761
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 9769 10795 9827 10801
rect 9769 10792 9781 10795
rect 7984 10764 9781 10792
rect 7984 10752 7990 10764
rect 9769 10761 9781 10764
rect 9815 10761 9827 10795
rect 10042 10792 10048 10804
rect 9769 10755 9827 10761
rect 9876 10764 10048 10792
rect 5092 10696 5212 10724
rect 5353 10727 5411 10733
rect 4801 10659 4859 10665
rect 4801 10625 4813 10659
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 4982 10616 4988 10668
rect 5040 10616 5046 10668
rect 5092 10665 5120 10696
rect 5353 10693 5365 10727
rect 5399 10724 5411 10727
rect 6270 10724 6276 10736
rect 5399 10696 6276 10724
rect 5399 10693 5411 10696
rect 5353 10687 5411 10693
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10625 5135 10659
rect 5077 10619 5135 10625
rect 5166 10616 5172 10668
rect 5224 10656 5230 10668
rect 5224 10628 5269 10656
rect 5224 10616 5230 10628
rect 3786 10588 3792 10600
rect 2792 10560 3792 10588
rect 3786 10548 3792 10560
rect 3844 10548 3850 10600
rect 3973 10591 4031 10597
rect 3973 10557 3985 10591
rect 4019 10588 4031 10591
rect 4540 10588 4568 10616
rect 4019 10560 4568 10588
rect 4617 10591 4675 10597
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 4617 10557 4629 10591
rect 4663 10588 4675 10591
rect 5368 10588 5396 10687
rect 6270 10684 6276 10696
rect 6328 10684 6334 10736
rect 8294 10724 8300 10736
rect 6840 10696 8300 10724
rect 5442 10616 5448 10668
rect 5500 10616 5506 10668
rect 5583 10659 5641 10665
rect 5583 10625 5595 10659
rect 5629 10656 5641 10659
rect 6086 10656 6092 10668
rect 5629 10628 6092 10656
rect 5629 10625 5641 10628
rect 5583 10619 5641 10625
rect 6086 10616 6092 10628
rect 6144 10656 6150 10668
rect 6840 10656 6868 10696
rect 8294 10684 8300 10696
rect 8352 10684 8358 10736
rect 9876 10724 9904 10764
rect 10042 10752 10048 10764
rect 10100 10752 10106 10804
rect 10870 10752 10876 10804
rect 10928 10792 10934 10804
rect 10928 10764 11652 10792
rect 10928 10752 10934 10764
rect 10594 10724 10600 10736
rect 8680 10696 8892 10724
rect 6144 10628 6868 10656
rect 6917 10659 6975 10665
rect 6144 10616 6150 10628
rect 6917 10625 6929 10659
rect 6963 10656 6975 10659
rect 7006 10656 7012 10668
rect 6963 10628 7012 10656
rect 6963 10625 6975 10628
rect 6917 10619 6975 10625
rect 7006 10616 7012 10628
rect 7064 10616 7070 10668
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10656 7159 10659
rect 8202 10656 8208 10668
rect 7147 10628 8208 10656
rect 7147 10625 7159 10628
rect 7101 10619 7159 10625
rect 8202 10616 8208 10628
rect 8260 10656 8266 10668
rect 8680 10656 8708 10696
rect 8260 10628 8708 10656
rect 8260 10616 8266 10628
rect 8754 10616 8760 10668
rect 8812 10616 8818 10668
rect 8864 10654 8892 10696
rect 9324 10696 9904 10724
rect 9963 10696 10600 10724
rect 8941 10659 8999 10665
rect 8941 10654 8953 10659
rect 8864 10626 8953 10654
rect 8941 10625 8953 10626
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 9214 10616 9220 10668
rect 9272 10616 9278 10668
rect 9324 10665 9352 10696
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10625 9367 10659
rect 9309 10619 9367 10625
rect 9398 10616 9404 10668
rect 9456 10616 9462 10668
rect 9963 10665 9991 10696
rect 10594 10684 10600 10696
rect 10652 10724 10658 10736
rect 11514 10724 11520 10736
rect 10652 10696 11520 10724
rect 10652 10684 10658 10696
rect 11514 10684 11520 10696
rect 11572 10684 11578 10736
rect 11624 10724 11652 10764
rect 11974 10752 11980 10804
rect 12032 10792 12038 10804
rect 12437 10795 12495 10801
rect 12437 10792 12449 10795
rect 12032 10764 12449 10792
rect 12032 10752 12038 10764
rect 12437 10761 12449 10764
rect 12483 10761 12495 10795
rect 12437 10755 12495 10761
rect 12529 10795 12587 10801
rect 12529 10761 12541 10795
rect 12575 10792 12587 10795
rect 12802 10792 12808 10804
rect 12575 10764 12808 10792
rect 12575 10761 12587 10764
rect 12529 10755 12587 10761
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 13740 10764 14412 10792
rect 11624 10696 12112 10724
rect 9948 10659 10006 10665
rect 9948 10625 9960 10659
rect 9994 10625 10006 10659
rect 9948 10619 10006 10625
rect 10042 10616 10048 10668
rect 10100 10616 10106 10668
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10625 10195 10659
rect 10137 10619 10195 10625
rect 4663 10560 5396 10588
rect 4663 10557 4675 10560
rect 4617 10551 4675 10557
rect 8570 10548 8576 10600
rect 8628 10588 8634 10600
rect 9125 10591 9183 10597
rect 9125 10588 9137 10591
rect 8628 10560 9137 10588
rect 8628 10548 8634 10560
rect 9125 10557 9137 10560
rect 9171 10588 9183 10591
rect 9490 10588 9496 10600
rect 9171 10560 9496 10588
rect 9171 10557 9183 10560
rect 9125 10551 9183 10557
rect 9490 10548 9496 10560
rect 9548 10548 9554 10600
rect 9582 10548 9588 10600
rect 9640 10548 9646 10600
rect 10152 10588 10180 10619
rect 10226 10616 10232 10668
rect 10284 10665 10290 10668
rect 10284 10659 10323 10665
rect 10311 10625 10323 10659
rect 10284 10619 10323 10625
rect 10413 10659 10471 10665
rect 10413 10625 10425 10659
rect 10459 10656 10471 10659
rect 10870 10656 10876 10668
rect 10459 10628 10876 10656
rect 10459 10625 10471 10628
rect 10413 10619 10471 10625
rect 10284 10616 10290 10619
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 10965 10659 11023 10665
rect 10965 10625 10977 10659
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 10060 10560 10180 10588
rect 4709 10523 4767 10529
rect 4709 10489 4721 10523
rect 4755 10520 4767 10523
rect 8938 10520 8944 10532
rect 4755 10492 8944 10520
rect 4755 10489 4767 10492
rect 4709 10483 4767 10489
rect 8938 10480 8944 10492
rect 8996 10480 9002 10532
rect 9600 10520 9628 10548
rect 10060 10520 10088 10560
rect 10686 10548 10692 10600
rect 10744 10588 10750 10600
rect 10980 10588 11008 10619
rect 11146 10616 11152 10668
rect 11204 10616 11210 10668
rect 11885 10659 11943 10665
rect 11885 10656 11897 10659
rect 11348 10628 11897 10656
rect 10744 10560 11008 10588
rect 10744 10548 10750 10560
rect 9143 10492 10088 10520
rect 3050 10412 3056 10464
rect 3108 10452 3114 10464
rect 3326 10452 3332 10464
rect 3108 10424 3332 10452
rect 3108 10412 3114 10424
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 3602 10412 3608 10464
rect 3660 10452 3666 10464
rect 3881 10455 3939 10461
rect 3881 10452 3893 10455
rect 3660 10424 3893 10452
rect 3660 10412 3666 10424
rect 3881 10421 3893 10424
rect 3927 10421 3939 10455
rect 3881 10415 3939 10421
rect 3970 10412 3976 10464
rect 4028 10452 4034 10464
rect 4249 10455 4307 10461
rect 4249 10452 4261 10455
rect 4028 10424 4261 10452
rect 4028 10412 4034 10424
rect 4249 10421 4261 10424
rect 4295 10421 4307 10455
rect 4249 10415 4307 10421
rect 4341 10455 4399 10461
rect 4341 10421 4353 10455
rect 4387 10452 4399 10455
rect 4798 10452 4804 10464
rect 4387 10424 4804 10452
rect 4387 10421 4399 10424
rect 4341 10415 4399 10421
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 6822 10412 6828 10464
rect 6880 10452 6886 10464
rect 8662 10452 8668 10464
rect 6880 10424 8668 10452
rect 6880 10412 6886 10424
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 8846 10412 8852 10464
rect 8904 10452 8910 10464
rect 9143 10452 9171 10492
rect 10134 10480 10140 10532
rect 10192 10520 10198 10532
rect 11348 10529 11376 10628
rect 11885 10625 11897 10628
rect 11931 10656 11943 10659
rect 11974 10656 11980 10668
rect 11931 10628 11980 10656
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 11974 10616 11980 10628
rect 12032 10616 12038 10668
rect 12084 10656 12112 10696
rect 12158 10684 12164 10736
rect 12216 10724 12222 10736
rect 12618 10724 12624 10736
rect 12216 10696 12624 10724
rect 12216 10684 12222 10696
rect 12618 10684 12624 10696
rect 12676 10733 12682 10736
rect 12676 10727 12739 10733
rect 12676 10693 12693 10727
rect 12727 10724 12739 10727
rect 12897 10727 12955 10733
rect 12727 10696 12769 10724
rect 12727 10693 12739 10696
rect 12676 10687 12739 10693
rect 12897 10693 12909 10727
rect 12943 10724 12955 10727
rect 13078 10724 13084 10736
rect 12943 10696 13084 10724
rect 12943 10693 12955 10696
rect 12897 10687 12955 10693
rect 12676 10684 12682 10687
rect 13078 10684 13084 10696
rect 13136 10684 13142 10736
rect 13740 10656 13768 10764
rect 13814 10684 13820 10736
rect 13872 10724 13878 10736
rect 14384 10724 14412 10764
rect 14918 10752 14924 10804
rect 14976 10792 14982 10804
rect 15289 10795 15347 10801
rect 15289 10792 15301 10795
rect 14976 10764 15301 10792
rect 14976 10752 14982 10764
rect 15289 10761 15301 10764
rect 15335 10761 15347 10795
rect 15289 10755 15347 10761
rect 15562 10752 15568 10804
rect 15620 10792 15626 10804
rect 16209 10795 16267 10801
rect 16209 10792 16221 10795
rect 15620 10764 16221 10792
rect 15620 10752 15626 10764
rect 16209 10761 16221 10764
rect 16255 10792 16267 10795
rect 17310 10792 17316 10804
rect 16255 10764 17316 10792
rect 16255 10761 16267 10764
rect 16209 10755 16267 10761
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 16945 10727 17003 10733
rect 13872 10696 14228 10724
rect 13872 10684 13878 10696
rect 12084 10628 13768 10656
rect 13998 10616 14004 10668
rect 14056 10616 14062 10668
rect 14200 10665 14228 10696
rect 14384 10696 15884 10724
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 14274 10616 14280 10668
rect 14332 10616 14338 10668
rect 14384 10665 14412 10696
rect 15304 10668 15332 10696
rect 14369 10659 14427 10665
rect 14369 10625 14381 10659
rect 14415 10625 14427 10659
rect 14369 10619 14427 10625
rect 15286 10616 15292 10668
rect 15344 10616 15350 10668
rect 15470 10616 15476 10668
rect 15528 10616 15534 10668
rect 15562 10616 15568 10668
rect 15620 10616 15626 10668
rect 15746 10616 15752 10668
rect 15804 10616 15810 10668
rect 15856 10665 15884 10696
rect 16945 10693 16957 10727
rect 16991 10724 17003 10727
rect 17126 10724 17132 10736
rect 16991 10696 17132 10724
rect 16991 10693 17003 10696
rect 16945 10687 17003 10693
rect 17126 10684 17132 10696
rect 17184 10724 17190 10736
rect 17402 10724 17408 10736
rect 17184 10696 17408 10724
rect 17184 10684 17190 10696
rect 17402 10684 17408 10696
rect 17460 10684 17466 10736
rect 15841 10659 15899 10665
rect 15841 10625 15853 10659
rect 15887 10625 15899 10659
rect 15841 10619 15899 10625
rect 16022 10616 16028 10668
rect 16080 10656 16086 10668
rect 16301 10659 16359 10665
rect 16301 10656 16313 10659
rect 16080 10628 16313 10656
rect 16080 10616 16086 10628
rect 16301 10625 16313 10628
rect 16347 10656 16359 10659
rect 16390 10656 16396 10668
rect 16347 10628 16396 10656
rect 16347 10625 16359 10628
rect 16301 10619 16359 10625
rect 16390 10616 16396 10628
rect 16448 10656 16454 10668
rect 17313 10659 17371 10665
rect 17313 10656 17325 10659
rect 16448 10628 17325 10656
rect 16448 10616 16454 10628
rect 17313 10625 17325 10628
rect 17359 10625 17371 10659
rect 17313 10619 17371 10625
rect 12066 10588 12072 10600
rect 11440 10560 12072 10588
rect 11333 10523 11391 10529
rect 10192 10492 11192 10520
rect 10192 10480 10198 10492
rect 8904 10424 9171 10452
rect 8904 10412 8910 10424
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 9585 10455 9643 10461
rect 9585 10452 9597 10455
rect 9272 10424 9597 10452
rect 9272 10412 9278 10424
rect 9585 10421 9597 10424
rect 9631 10421 9643 10455
rect 9585 10415 9643 10421
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 10686 10452 10692 10464
rect 9824 10424 10692 10452
rect 9824 10412 9830 10424
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 11054 10412 11060 10464
rect 11112 10412 11118 10464
rect 11164 10452 11192 10492
rect 11333 10489 11345 10523
rect 11379 10489 11391 10523
rect 11333 10483 11391 10489
rect 11440 10452 11468 10560
rect 12066 10548 12072 10560
rect 12124 10548 12130 10600
rect 12161 10591 12219 10597
rect 12161 10557 12173 10591
rect 12207 10588 12219 10591
rect 15194 10588 15200 10600
rect 12207 10560 15200 10588
rect 12207 10557 12219 10560
rect 12161 10551 12219 10557
rect 15194 10548 15200 10560
rect 15252 10588 15258 10600
rect 16828 10591 16886 10597
rect 15252 10560 16712 10588
rect 15252 10548 15258 10560
rect 16114 10520 16120 10532
rect 12268 10492 16120 10520
rect 11164 10424 11468 10452
rect 11790 10412 11796 10464
rect 11848 10452 11854 10464
rect 12268 10461 12296 10492
rect 16114 10480 16120 10492
rect 16172 10480 16178 10532
rect 16684 10529 16712 10560
rect 16828 10557 16840 10591
rect 16874 10557 16886 10591
rect 16828 10551 16886 10557
rect 16669 10523 16727 10529
rect 16669 10489 16681 10523
rect 16715 10489 16727 10523
rect 16843 10520 16871 10551
rect 17034 10548 17040 10600
rect 17092 10548 17098 10600
rect 17586 10520 17592 10532
rect 16843 10492 17592 10520
rect 16669 10483 16727 10489
rect 17586 10480 17592 10492
rect 17644 10480 17650 10532
rect 12253 10455 12311 10461
rect 12253 10452 12265 10455
rect 11848 10424 12265 10452
rect 11848 10412 11854 10424
rect 12253 10421 12265 10424
rect 12299 10421 12311 10455
rect 12253 10415 12311 10421
rect 12710 10412 12716 10464
rect 12768 10412 12774 10464
rect 12894 10412 12900 10464
rect 12952 10452 12958 10464
rect 13630 10452 13636 10464
rect 12952 10424 13636 10452
rect 12952 10412 12958 10424
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 14090 10412 14096 10464
rect 14148 10452 14154 10464
rect 14645 10455 14703 10461
rect 14645 10452 14657 10455
rect 14148 10424 14657 10452
rect 14148 10412 14154 10424
rect 14645 10421 14657 10424
rect 14691 10421 14703 10455
rect 14645 10415 14703 10421
rect 14734 10412 14740 10464
rect 14792 10452 14798 10464
rect 17126 10452 17132 10464
rect 14792 10424 17132 10452
rect 14792 10412 14798 10424
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 1104 10362 18400 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 18400 10362
rect 1104 10288 18400 10310
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 3329 10251 3387 10257
rect 3329 10248 3341 10251
rect 2832 10220 3341 10248
rect 2832 10208 2838 10220
rect 3329 10217 3341 10220
rect 3375 10217 3387 10251
rect 3329 10211 3387 10217
rect 4246 10208 4252 10260
rect 4304 10248 4310 10260
rect 4798 10248 4804 10260
rect 4304 10220 4804 10248
rect 4304 10208 4310 10220
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 6178 10208 6184 10260
rect 6236 10248 6242 10260
rect 6822 10248 6828 10260
rect 6236 10220 6828 10248
rect 6236 10208 6242 10220
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 7282 10248 7288 10260
rect 6972 10220 7288 10248
rect 6972 10208 6978 10220
rect 7282 10208 7288 10220
rect 7340 10248 7346 10260
rect 7469 10251 7527 10257
rect 7469 10248 7481 10251
rect 7340 10220 7481 10248
rect 7340 10208 7346 10220
rect 7469 10217 7481 10220
rect 7515 10217 7527 10251
rect 7469 10211 7527 10217
rect 7926 10208 7932 10260
rect 7984 10248 7990 10260
rect 7984 10220 9352 10248
rect 7984 10208 7990 10220
rect 3970 10140 3976 10192
rect 4028 10140 4034 10192
rect 5718 10180 5724 10192
rect 4172 10152 5724 10180
rect 2406 10072 2412 10124
rect 2464 10112 2470 10124
rect 2685 10115 2743 10121
rect 2685 10112 2697 10115
rect 2464 10084 2697 10112
rect 2464 10072 2470 10084
rect 2685 10081 2697 10084
rect 2731 10081 2743 10115
rect 2685 10075 2743 10081
rect 2823 10115 2881 10121
rect 2823 10081 2835 10115
rect 2869 10112 2881 10115
rect 3510 10112 3516 10124
rect 2869 10084 3516 10112
rect 2869 10081 2881 10084
rect 2823 10075 2881 10081
rect 3510 10072 3516 10084
rect 3568 10072 3574 10124
rect 3988 10112 4016 10140
rect 4172 10121 4200 10152
rect 5718 10140 5724 10152
rect 5776 10140 5782 10192
rect 5994 10140 6000 10192
rect 6052 10180 6058 10192
rect 6270 10180 6276 10192
rect 6052 10152 6276 10180
rect 6052 10140 6058 10152
rect 6270 10140 6276 10152
rect 6328 10140 6334 10192
rect 8570 10180 8576 10192
rect 7024 10152 8576 10180
rect 4065 10115 4123 10121
rect 4065 10112 4077 10115
rect 3988 10084 4077 10112
rect 4065 10081 4077 10084
rect 4111 10081 4123 10115
rect 4065 10075 4123 10081
rect 4157 10115 4215 10121
rect 4157 10081 4169 10115
rect 4203 10081 4215 10115
rect 4157 10075 4215 10081
rect 4246 10072 4252 10124
rect 4304 10072 4310 10124
rect 4706 10072 4712 10124
rect 4764 10112 4770 10124
rect 4764 10084 5028 10112
rect 4764 10072 4770 10084
rect 2501 10047 2559 10053
rect 2501 10013 2513 10047
rect 2547 10013 2559 10047
rect 2501 10007 2559 10013
rect 2516 9976 2544 10007
rect 2958 10004 2964 10056
rect 3016 10004 3022 10056
rect 3050 10004 3056 10056
rect 3108 10004 3114 10056
rect 3326 10004 3332 10056
rect 3384 10004 3390 10056
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10013 4031 10047
rect 3973 10007 4031 10013
rect 3145 9979 3203 9985
rect 3145 9976 3157 9979
rect 2516 9948 3157 9976
rect 3145 9945 3157 9948
rect 3191 9976 3203 9979
rect 3878 9976 3884 9988
rect 3191 9948 3884 9976
rect 3191 9945 3203 9948
rect 3145 9939 3203 9945
rect 3878 9936 3884 9948
rect 3936 9936 3942 9988
rect 3988 9976 4016 10007
rect 4430 10004 4436 10056
rect 4488 10044 4494 10056
rect 4798 10053 4804 10056
rect 4617 10047 4675 10053
rect 4617 10044 4629 10047
rect 4488 10016 4629 10044
rect 4488 10004 4494 10016
rect 4617 10013 4629 10016
rect 4663 10013 4675 10047
rect 4796 10044 4804 10053
rect 4617 10007 4675 10013
rect 4724 10016 4804 10044
rect 4246 9976 4252 9988
rect 3988 9948 4252 9976
rect 4246 9936 4252 9948
rect 4304 9936 4310 9988
rect 4724 9976 4752 10016
rect 4796 10007 4804 10016
rect 4798 10004 4804 10007
rect 4856 10004 4862 10056
rect 4890 10004 4896 10056
rect 4948 10004 4954 10056
rect 5000 10053 5028 10084
rect 5442 10072 5448 10124
rect 5500 10112 5506 10124
rect 5810 10112 5816 10124
rect 5500 10084 5816 10112
rect 5500 10072 5506 10084
rect 5810 10072 5816 10084
rect 5868 10112 5874 10124
rect 6917 10115 6975 10121
rect 6917 10112 6929 10115
rect 5868 10084 6929 10112
rect 5868 10072 5874 10084
rect 6917 10081 6929 10084
rect 6963 10081 6975 10115
rect 6917 10075 6975 10081
rect 7024 10053 7052 10152
rect 8570 10140 8576 10152
rect 8628 10140 8634 10192
rect 9122 10140 9128 10192
rect 9180 10180 9186 10192
rect 9217 10183 9275 10189
rect 9217 10180 9229 10183
rect 9180 10152 9229 10180
rect 9180 10140 9186 10152
rect 9217 10149 9229 10152
rect 9263 10149 9275 10183
rect 9324 10180 9352 10220
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 9677 10251 9735 10257
rect 9677 10248 9689 10251
rect 9548 10220 9689 10248
rect 9548 10208 9554 10220
rect 9677 10217 9689 10220
rect 9723 10217 9735 10251
rect 9677 10211 9735 10217
rect 10594 10208 10600 10260
rect 10652 10248 10658 10260
rect 10652 10220 13216 10248
rect 10652 10208 10658 10220
rect 13188 10192 13216 10220
rect 14550 10208 14556 10260
rect 14608 10208 14614 10260
rect 15746 10208 15752 10260
rect 15804 10248 15810 10260
rect 16206 10248 16212 10260
rect 15804 10220 16212 10248
rect 15804 10208 15810 10220
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 16298 10208 16304 10260
rect 16356 10248 16362 10260
rect 16393 10251 16451 10257
rect 16393 10248 16405 10251
rect 16356 10220 16405 10248
rect 16356 10208 16362 10220
rect 16393 10217 16405 10220
rect 16439 10217 16451 10251
rect 16393 10211 16451 10217
rect 9858 10180 9864 10192
rect 9324 10152 9864 10180
rect 9217 10143 9275 10149
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 10870 10180 10876 10192
rect 9968 10152 10876 10180
rect 8665 10115 8723 10121
rect 8665 10081 8677 10115
rect 8711 10112 8723 10115
rect 9309 10115 9367 10121
rect 9309 10112 9321 10115
rect 8711 10084 9321 10112
rect 8711 10081 8723 10084
rect 8665 10075 8723 10081
rect 9309 10081 9321 10084
rect 9355 10081 9367 10115
rect 9968 10112 9996 10152
rect 10870 10140 10876 10152
rect 10928 10140 10934 10192
rect 11164 10152 12388 10180
rect 9309 10075 9367 10081
rect 9416 10084 9996 10112
rect 9416 10056 9444 10084
rect 10042 10072 10048 10124
rect 10100 10072 10106 10124
rect 11164 10121 11192 10152
rect 11149 10115 11207 10121
rect 11149 10081 11161 10115
rect 11195 10081 11207 10115
rect 11149 10075 11207 10081
rect 11241 10115 11299 10121
rect 11241 10081 11253 10115
rect 11287 10112 11299 10115
rect 11514 10112 11520 10124
rect 11287 10084 11520 10112
rect 11287 10081 11299 10084
rect 11241 10075 11299 10081
rect 11514 10072 11520 10084
rect 11572 10072 11578 10124
rect 11609 10115 11667 10121
rect 11609 10081 11621 10115
rect 11655 10112 11667 10115
rect 12360 10112 12388 10152
rect 13170 10140 13176 10192
rect 13228 10140 13234 10192
rect 14568 10180 14596 10208
rect 16761 10183 16819 10189
rect 16761 10180 16773 10183
rect 14568 10152 16773 10180
rect 16761 10149 16773 10152
rect 16807 10180 16819 10183
rect 17034 10180 17040 10192
rect 16807 10152 17040 10180
rect 16807 10149 16819 10152
rect 16761 10143 16819 10149
rect 17034 10140 17040 10152
rect 17092 10140 17098 10192
rect 12986 10112 12992 10124
rect 11655 10084 12296 10112
rect 12360 10084 12992 10112
rect 11655 10081 11667 10084
rect 11609 10075 11667 10081
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10013 5043 10047
rect 7009 10047 7067 10053
rect 4985 10007 5043 10013
rect 5092 10016 6960 10044
rect 5092 9976 5120 10016
rect 4724 9948 5120 9976
rect 5626 9936 5632 9988
rect 5684 9976 5690 9988
rect 5721 9979 5779 9985
rect 5721 9976 5733 9979
rect 5684 9948 5733 9976
rect 5684 9936 5690 9948
rect 5721 9945 5733 9948
rect 5767 9945 5779 9979
rect 5721 9939 5779 9945
rect 6273 9979 6331 9985
rect 6273 9945 6285 9979
rect 6319 9976 6331 9979
rect 6822 9976 6828 9988
rect 6319 9948 6828 9976
rect 6319 9945 6331 9948
rect 6273 9939 6331 9945
rect 6822 9936 6828 9948
rect 6880 9936 6886 9988
rect 6932 9976 6960 10016
rect 7009 10013 7021 10047
rect 7055 10013 7067 10047
rect 7009 10007 7067 10013
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10044 7159 10047
rect 7190 10044 7196 10056
rect 7147 10016 7196 10044
rect 7147 10013 7159 10016
rect 7101 10007 7159 10013
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 7282 10004 7288 10056
rect 7340 10004 7346 10056
rect 8570 10044 8576 10056
rect 7392 10016 8576 10044
rect 7392 9976 7420 10016
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 8754 10004 8760 10056
rect 8812 10004 8818 10056
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 6932 9948 7420 9976
rect 7558 9936 7564 9988
rect 7616 9936 7622 9988
rect 7742 9936 7748 9988
rect 7800 9976 7806 9988
rect 8956 9976 8984 10007
rect 9030 10004 9036 10056
rect 9088 10044 9094 10056
rect 9125 10047 9183 10053
rect 9125 10044 9137 10047
rect 9088 10016 9137 10044
rect 9088 10004 9094 10016
rect 9125 10013 9137 10016
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 9398 10004 9404 10056
rect 9456 10004 9462 10056
rect 9490 10004 9496 10056
rect 9548 10044 9554 10056
rect 10060 10044 10088 10072
rect 9548 10016 10088 10044
rect 10873 10047 10931 10053
rect 9548 10004 9554 10016
rect 10873 10013 10885 10047
rect 10919 10013 10931 10047
rect 10873 10007 10931 10013
rect 7800 9948 8984 9976
rect 7800 9936 7806 9948
rect 2498 9868 2504 9920
rect 2556 9868 2562 9920
rect 3694 9868 3700 9920
rect 3752 9908 3758 9920
rect 3789 9911 3847 9917
rect 3789 9908 3801 9911
rect 3752 9880 3801 9908
rect 3752 9868 3758 9880
rect 3789 9877 3801 9880
rect 3835 9877 3847 9911
rect 3789 9871 3847 9877
rect 4706 9868 4712 9920
rect 4764 9908 4770 9920
rect 4890 9908 4896 9920
rect 4764 9880 4896 9908
rect 4764 9868 4770 9880
rect 4890 9868 4896 9880
rect 4948 9868 4954 9920
rect 5258 9868 5264 9920
rect 5316 9868 5322 9920
rect 5445 9911 5503 9917
rect 5445 9877 5457 9911
rect 5491 9908 5503 9911
rect 5534 9908 5540 9920
rect 5491 9880 5540 9908
rect 5491 9877 5503 9880
rect 5445 9871 5503 9877
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 5994 9868 6000 9920
rect 6052 9868 6058 9920
rect 6546 9868 6552 9920
rect 6604 9908 6610 9920
rect 6641 9911 6699 9917
rect 6641 9908 6653 9911
rect 6604 9880 6653 9908
rect 6604 9868 6610 9880
rect 6641 9877 6653 9880
rect 6687 9877 6699 9911
rect 6641 9871 6699 9877
rect 7006 9868 7012 9920
rect 7064 9908 7070 9920
rect 7190 9908 7196 9920
rect 7064 9880 7196 9908
rect 7064 9868 7070 9880
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 7282 9868 7288 9920
rect 7340 9868 7346 9920
rect 8956 9908 8984 9948
rect 9674 9936 9680 9988
rect 9732 9976 9738 9988
rect 9953 9979 10011 9985
rect 9953 9976 9965 9979
rect 9732 9948 9965 9976
rect 9732 9936 9738 9948
rect 9953 9945 9965 9948
rect 9999 9976 10011 9979
rect 10888 9976 10916 10007
rect 11054 10004 11060 10056
rect 11112 10004 11118 10056
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 11425 10047 11483 10053
rect 11425 10044 11437 10047
rect 11388 10016 11437 10044
rect 11388 10004 11394 10016
rect 11425 10013 11437 10016
rect 11471 10044 11483 10047
rect 11698 10044 11704 10056
rect 11471 10016 11704 10044
rect 11471 10013 11483 10016
rect 11425 10007 11483 10013
rect 11698 10004 11704 10016
rect 11756 10004 11762 10056
rect 11882 10004 11888 10056
rect 11940 10004 11946 10056
rect 11974 10004 11980 10056
rect 12032 10004 12038 10056
rect 12268 10053 12296 10084
rect 12253 10047 12311 10053
rect 12253 10013 12265 10047
rect 12299 10013 12311 10047
rect 12253 10007 12311 10013
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10013 12403 10047
rect 12345 10007 12403 10013
rect 11790 9976 11796 9988
rect 9999 9948 11796 9976
rect 9999 9945 10011 9948
rect 9953 9939 10011 9945
rect 11790 9936 11796 9948
rect 11848 9936 11854 9988
rect 12066 9936 12072 9988
rect 12124 9936 12130 9988
rect 12158 9936 12164 9988
rect 12216 9976 12222 9988
rect 12360 9976 12388 10007
rect 12618 10004 12624 10056
rect 12676 10004 12682 10056
rect 12820 10053 12848 10084
rect 12986 10072 12992 10084
rect 13044 10072 13050 10124
rect 13998 10112 14004 10124
rect 13464 10084 14004 10112
rect 12805 10047 12863 10053
rect 12805 10013 12817 10047
rect 12851 10013 12863 10047
rect 12805 10007 12863 10013
rect 13078 10004 13084 10056
rect 13136 10004 13142 10056
rect 13464 10053 13492 10084
rect 13998 10072 14004 10084
rect 14056 10112 14062 10124
rect 14550 10112 14556 10124
rect 14056 10084 14556 10112
rect 14056 10072 14062 10084
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 14660 10084 15424 10112
rect 13448 10047 13506 10053
rect 13448 10013 13460 10047
rect 13494 10013 13506 10047
rect 13448 10007 13506 10013
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10044 13599 10047
rect 13630 10044 13636 10056
rect 13587 10016 13636 10044
rect 13587 10013 13599 10016
rect 13541 10007 13599 10013
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 14660 10053 14688 10084
rect 15396 10056 15424 10084
rect 14644 10047 14702 10053
rect 14644 10013 14656 10047
rect 14690 10013 14702 10047
rect 14644 10007 14702 10013
rect 14734 10004 14740 10056
rect 14792 10004 14798 10056
rect 15378 10004 15384 10056
rect 15436 10004 15442 10056
rect 15470 10004 15476 10056
rect 15528 10044 15534 10056
rect 15565 10047 15623 10053
rect 15565 10044 15577 10047
rect 15528 10016 15577 10044
rect 15528 10004 15534 10016
rect 15565 10013 15577 10016
rect 15611 10013 15623 10047
rect 15565 10007 15623 10013
rect 15838 10004 15844 10056
rect 15896 10044 15902 10056
rect 15933 10047 15991 10053
rect 15933 10044 15945 10047
rect 15896 10016 15945 10044
rect 15896 10004 15902 10016
rect 15933 10013 15945 10016
rect 15979 10044 15991 10047
rect 16853 10047 16911 10053
rect 16853 10044 16865 10047
rect 15979 10016 16865 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 16853 10013 16865 10016
rect 16899 10013 16911 10047
rect 16853 10007 16911 10013
rect 17218 10004 17224 10056
rect 17276 10004 17282 10056
rect 12216 9948 12388 9976
rect 12713 9979 12771 9985
rect 12216 9936 12222 9948
rect 12713 9945 12725 9979
rect 12759 9945 12771 9979
rect 12713 9939 12771 9945
rect 12943 9979 13001 9985
rect 12943 9945 12955 9979
rect 12989 9976 13001 9979
rect 14366 9976 14372 9988
rect 12989 9948 14372 9976
rect 12989 9945 13001 9948
rect 12943 9939 13001 9945
rect 9861 9911 9919 9917
rect 9861 9908 9873 9911
rect 8956 9880 9873 9908
rect 9861 9877 9873 9880
rect 9907 9877 9919 9911
rect 9861 9871 9919 9877
rect 10226 9868 10232 9920
rect 10284 9908 10290 9920
rect 11701 9911 11759 9917
rect 11701 9908 11713 9911
rect 10284 9880 11713 9908
rect 10284 9868 10290 9880
rect 11701 9877 11713 9880
rect 11747 9877 11759 9911
rect 11701 9871 11759 9877
rect 12434 9868 12440 9920
rect 12492 9868 12498 9920
rect 12728 9908 12756 9939
rect 14366 9936 14372 9948
rect 14424 9936 14430 9988
rect 15194 9936 15200 9988
rect 15252 9976 15258 9988
rect 15289 9979 15347 9985
rect 15289 9976 15301 9979
rect 15252 9948 15301 9976
rect 15252 9936 15258 9948
rect 15289 9945 15301 9948
rect 15335 9945 15347 9979
rect 15289 9939 15347 9945
rect 16390 9936 16396 9988
rect 16448 9976 16454 9988
rect 16942 9976 16948 9988
rect 16448 9948 16948 9976
rect 16448 9936 16454 9948
rect 16942 9936 16948 9948
rect 17000 9936 17006 9988
rect 13173 9911 13231 9917
rect 13173 9908 13185 9911
rect 12728 9880 13185 9908
rect 13173 9877 13185 9880
rect 13219 9877 13231 9911
rect 13173 9871 13231 9877
rect 16022 9868 16028 9920
rect 16080 9868 16086 9920
rect 1104 9818 18400 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 18400 9818
rect 1104 9744 18400 9766
rect 2961 9707 3019 9713
rect 2961 9673 2973 9707
rect 3007 9704 3019 9707
rect 3050 9704 3056 9716
rect 3007 9676 3056 9704
rect 3007 9673 3019 9676
rect 2961 9667 3019 9673
rect 3050 9664 3056 9676
rect 3108 9664 3114 9716
rect 3602 9664 3608 9716
rect 3660 9704 3666 9716
rect 3789 9707 3847 9713
rect 3789 9704 3801 9707
rect 3660 9676 3801 9704
rect 3660 9664 3666 9676
rect 3789 9673 3801 9676
rect 3835 9673 3847 9707
rect 3789 9667 3847 9673
rect 4614 9664 4620 9716
rect 4672 9704 4678 9716
rect 4890 9704 4896 9716
rect 4672 9676 4896 9704
rect 4672 9664 4678 9676
rect 4890 9664 4896 9676
rect 4948 9704 4954 9716
rect 6454 9704 6460 9716
rect 4948 9676 6460 9704
rect 4948 9664 4954 9676
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 6822 9664 6828 9716
rect 6880 9704 6886 9716
rect 7926 9704 7932 9716
rect 6880 9676 7932 9704
rect 6880 9664 6886 9676
rect 7926 9664 7932 9676
rect 7984 9664 7990 9716
rect 9582 9664 9588 9716
rect 9640 9704 9646 9716
rect 9861 9707 9919 9713
rect 9861 9704 9873 9707
rect 9640 9676 9873 9704
rect 9640 9664 9646 9676
rect 9861 9673 9873 9676
rect 9907 9673 9919 9707
rect 9861 9667 9919 9673
rect 11514 9664 11520 9716
rect 11572 9704 11578 9716
rect 11974 9704 11980 9716
rect 11572 9676 11980 9704
rect 11572 9664 11578 9676
rect 11974 9664 11980 9676
rect 12032 9664 12038 9716
rect 12618 9704 12624 9716
rect 12360 9676 12624 9704
rect 2317 9639 2375 9645
rect 2317 9636 2329 9639
rect 1688 9608 2329 9636
rect 1688 9577 1716 9608
rect 2317 9605 2329 9608
rect 2363 9605 2375 9639
rect 3694 9636 3700 9648
rect 2317 9599 2375 9605
rect 2424 9608 2636 9636
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9537 1731 9571
rect 1673 9531 1731 9537
rect 2222 9528 2228 9580
rect 2280 9568 2286 9580
rect 2424 9568 2452 9608
rect 2280 9540 2452 9568
rect 2280 9528 2286 9540
rect 2498 9528 2504 9580
rect 2556 9528 2562 9580
rect 2608 9577 2636 9608
rect 2884 9608 3700 9636
rect 2884 9580 2912 9608
rect 3694 9596 3700 9608
rect 3752 9596 3758 9648
rect 4246 9596 4252 9648
rect 4304 9596 4310 9648
rect 5445 9639 5503 9645
rect 5445 9636 5457 9639
rect 4448 9608 5457 9636
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9537 2651 9571
rect 2593 9531 2651 9537
rect 2682 9528 2688 9580
rect 2740 9568 2746 9580
rect 2777 9571 2835 9577
rect 2777 9568 2789 9571
rect 2740 9540 2789 9568
rect 2740 9528 2746 9540
rect 2777 9537 2789 9540
rect 2823 9537 2835 9571
rect 2777 9531 2835 9537
rect 2866 9528 2872 9580
rect 2924 9528 2930 9580
rect 3050 9528 3056 9580
rect 3108 9568 3114 9580
rect 3145 9571 3203 9577
rect 3145 9568 3157 9571
rect 3108 9540 3157 9568
rect 3108 9528 3114 9540
rect 3145 9537 3157 9540
rect 3191 9537 3203 9571
rect 3145 9531 3203 9537
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9568 3295 9571
rect 3326 9568 3332 9580
rect 3283 9540 3332 9568
rect 3283 9537 3295 9540
rect 3237 9531 3295 9537
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 3513 9571 3571 9577
rect 3513 9537 3525 9571
rect 3559 9537 3571 9571
rect 3513 9531 3571 9537
rect 1762 9460 1768 9512
rect 1820 9460 1826 9512
rect 2133 9503 2191 9509
rect 2133 9469 2145 9503
rect 2179 9500 2191 9503
rect 2314 9500 2320 9512
rect 2179 9472 2320 9500
rect 2179 9469 2191 9472
rect 2133 9463 2191 9469
rect 2314 9460 2320 9472
rect 2372 9460 2378 9512
rect 2406 9460 2412 9512
rect 2464 9500 2470 9512
rect 3436 9500 3464 9531
rect 2464 9472 3464 9500
rect 2464 9460 2470 9472
rect 2958 9392 2964 9444
rect 3016 9432 3022 9444
rect 3528 9432 3556 9531
rect 3602 9528 3608 9580
rect 3660 9528 3666 9580
rect 4448 9577 4476 9608
rect 5445 9605 5457 9608
rect 5491 9605 5503 9639
rect 5445 9599 5503 9605
rect 5810 9596 5816 9648
rect 5868 9596 5874 9648
rect 7837 9639 7895 9645
rect 7837 9636 7849 9639
rect 7208 9608 7849 9636
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 4614 9528 4620 9580
rect 4672 9528 4678 9580
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 5166 9568 5172 9580
rect 4755 9540 5172 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9537 5319 9571
rect 5629 9571 5687 9577
rect 5629 9568 5641 9571
rect 5261 9531 5319 9537
rect 5552 9540 5641 9568
rect 4798 9460 4804 9512
rect 4856 9500 4862 9512
rect 4893 9503 4951 9509
rect 4893 9500 4905 9503
rect 4856 9472 4905 9500
rect 4856 9460 4862 9472
rect 4893 9469 4905 9472
rect 4939 9469 4951 9503
rect 4893 9463 4951 9469
rect 4982 9460 4988 9512
rect 5040 9460 5046 9512
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 5276 9500 5304 9531
rect 5132 9472 5304 9500
rect 5132 9460 5138 9472
rect 3970 9432 3976 9444
rect 3016 9404 3976 9432
rect 3016 9392 3022 9404
rect 3970 9392 3976 9404
rect 4028 9432 4034 9444
rect 5552 9432 5580 9540
rect 5629 9537 5641 9540
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 5902 9528 5908 9580
rect 5960 9528 5966 9580
rect 6454 9528 6460 9580
rect 6512 9568 6518 9580
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6512 9540 6561 9568
rect 6512 9528 6518 9540
rect 6549 9537 6561 9540
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 7006 9568 7012 9580
rect 6687 9540 7012 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 7208 9568 7236 9608
rect 7837 9605 7849 9608
rect 7883 9636 7895 9639
rect 12360 9636 12388 9676
rect 12618 9664 12624 9676
rect 12676 9704 12682 9716
rect 13078 9704 13084 9716
rect 12676 9676 13084 9704
rect 12676 9664 12682 9676
rect 13078 9664 13084 9676
rect 13136 9664 13142 9716
rect 13354 9664 13360 9716
rect 13412 9704 13418 9716
rect 14458 9704 14464 9716
rect 13412 9676 14464 9704
rect 13412 9664 13418 9676
rect 7883 9608 12388 9636
rect 7883 9605 7895 9608
rect 7837 9599 7895 9605
rect 12434 9596 12440 9648
rect 12492 9596 12498 9648
rect 12526 9596 12532 9648
rect 12584 9596 12590 9648
rect 7117 9540 7236 9568
rect 6733 9503 6791 9509
rect 6733 9469 6745 9503
rect 6779 9469 6791 9503
rect 6733 9463 6791 9469
rect 6748 9432 6776 9463
rect 6822 9460 6828 9512
rect 6880 9460 6886 9512
rect 7117 9500 7145 9540
rect 7282 9528 7288 9580
rect 7340 9528 7346 9580
rect 7558 9528 7564 9580
rect 7616 9528 7622 9580
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9568 7803 9571
rect 7926 9568 7932 9580
rect 7791 9540 7932 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 9674 9528 9680 9580
rect 9732 9568 9738 9580
rect 9769 9571 9827 9577
rect 9769 9568 9781 9571
rect 9732 9540 9781 9568
rect 9732 9528 9738 9540
rect 9769 9537 9781 9540
rect 9815 9568 9827 9571
rect 10042 9568 10048 9580
rect 9815 9540 10048 9568
rect 9815 9537 9827 9540
rect 9769 9531 9827 9537
rect 10042 9528 10048 9540
rect 10100 9528 10106 9580
rect 10137 9571 10195 9577
rect 10137 9537 10149 9571
rect 10183 9568 10195 9571
rect 10962 9568 10968 9580
rect 10183 9540 10968 9568
rect 10183 9537 10195 9540
rect 10137 9531 10195 9537
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 12066 9528 12072 9580
rect 12124 9568 12130 9580
rect 12250 9568 12256 9580
rect 12124 9540 12256 9568
rect 12124 9528 12130 9540
rect 12250 9528 12256 9540
rect 12308 9528 12314 9580
rect 12621 9571 12679 9577
rect 12621 9537 12633 9571
rect 12667 9537 12679 9571
rect 12621 9531 12679 9537
rect 13173 9571 13231 9577
rect 13173 9537 13185 9571
rect 13219 9568 13231 9571
rect 13354 9568 13360 9580
rect 13219 9540 13360 9568
rect 13219 9537 13231 9540
rect 13173 9531 13231 9537
rect 6932 9472 7145 9500
rect 7193 9503 7251 9509
rect 6932 9432 6960 9472
rect 7193 9469 7205 9503
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 4028 9404 6592 9432
rect 6748 9404 6960 9432
rect 4028 9392 4034 9404
rect 1489 9367 1547 9373
rect 1489 9333 1501 9367
rect 1535 9364 1547 9367
rect 1670 9364 1676 9376
rect 1535 9336 1676 9364
rect 1535 9333 1547 9336
rect 1489 9327 1547 9333
rect 1670 9324 1676 9336
rect 1728 9324 1734 9376
rect 3326 9324 3332 9376
rect 3384 9364 3390 9376
rect 3510 9364 3516 9376
rect 3384 9336 3516 9364
rect 3384 9324 3390 9336
rect 3510 9324 3516 9336
rect 3568 9364 3574 9376
rect 4982 9364 4988 9376
rect 3568 9336 4988 9364
rect 3568 9324 3574 9336
rect 4982 9324 4988 9336
rect 5040 9364 5046 9376
rect 5534 9364 5540 9376
rect 5040 9336 5540 9364
rect 5040 9324 5046 9336
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 6365 9367 6423 9373
rect 6365 9333 6377 9367
rect 6411 9364 6423 9367
rect 6454 9364 6460 9376
rect 6411 9336 6460 9364
rect 6411 9333 6423 9336
rect 6365 9327 6423 9333
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 6564 9364 6592 9404
rect 7006 9392 7012 9444
rect 7064 9392 7070 9444
rect 7208 9432 7236 9463
rect 7650 9460 7656 9512
rect 7708 9460 7714 9512
rect 9953 9503 10011 9509
rect 9953 9469 9965 9503
rect 9999 9500 10011 9503
rect 10778 9500 10784 9512
rect 9999 9472 10784 9500
rect 9999 9469 10011 9472
rect 9953 9463 10011 9469
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 11698 9460 11704 9512
rect 11756 9500 11762 9512
rect 12526 9500 12532 9512
rect 11756 9472 12532 9500
rect 11756 9460 11762 9472
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 12636 9500 12664 9531
rect 13354 9528 13360 9540
rect 13412 9528 13418 9580
rect 13998 9577 14004 9586
rect 13901 9571 13959 9577
rect 13901 9537 13913 9571
rect 13947 9537 13959 9571
rect 13901 9531 13959 9537
rect 13993 9534 14004 9577
rect 14056 9534 14062 9586
rect 14108 9568 14136 9676
rect 14458 9664 14464 9676
rect 14516 9664 14522 9716
rect 14550 9664 14556 9716
rect 14608 9704 14614 9716
rect 14921 9707 14979 9713
rect 14921 9704 14933 9707
rect 14608 9676 14933 9704
rect 14608 9664 14614 9676
rect 14921 9673 14933 9676
rect 14967 9673 14979 9707
rect 14921 9667 14979 9673
rect 16114 9596 16120 9648
rect 16172 9596 16178 9648
rect 14185 9571 14243 9577
rect 14185 9568 14197 9571
rect 14108 9540 14197 9568
rect 14185 9537 14197 9540
rect 14231 9537 14243 9571
rect 13993 9531 14051 9534
rect 14185 9531 14243 9537
rect 12710 9500 12716 9512
rect 12636 9472 12716 9500
rect 12710 9460 12716 9472
rect 12768 9500 12774 9512
rect 13924 9500 13952 9531
rect 14274 9528 14280 9580
rect 14332 9528 14338 9580
rect 14366 9528 14372 9580
rect 14424 9528 14430 9580
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9568 14519 9571
rect 14550 9568 14556 9580
rect 14507 9540 14556 9568
rect 14507 9537 14519 9540
rect 14461 9531 14519 9537
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 14642 9528 14648 9580
rect 14700 9528 14706 9580
rect 14734 9528 14740 9580
rect 14792 9528 14798 9580
rect 14918 9528 14924 9580
rect 14976 9568 14982 9580
rect 14976 9540 15700 9568
rect 14976 9528 14982 9540
rect 15010 9500 15016 9512
rect 12768 9472 13860 9500
rect 13924 9472 15016 9500
rect 12768 9460 12774 9472
rect 9030 9432 9036 9444
rect 7208 9404 9036 9432
rect 9030 9392 9036 9404
rect 9088 9392 9094 9444
rect 9858 9392 9864 9444
rect 9916 9432 9922 9444
rect 12989 9435 13047 9441
rect 9916 9404 12480 9432
rect 9916 9392 9922 9404
rect 6822 9364 6828 9376
rect 6564 9336 6828 9364
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 7374 9324 7380 9376
rect 7432 9364 7438 9376
rect 8110 9364 8116 9376
rect 7432 9336 8116 9364
rect 7432 9324 7438 9336
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 10042 9324 10048 9376
rect 10100 9364 10106 9376
rect 10137 9367 10195 9373
rect 10137 9364 10149 9367
rect 10100 9336 10149 9364
rect 10100 9324 10106 9336
rect 10137 9333 10149 9336
rect 10183 9333 10195 9367
rect 10137 9327 10195 9333
rect 11054 9324 11060 9376
rect 11112 9364 11118 9376
rect 11606 9364 11612 9376
rect 11112 9336 11612 9364
rect 11112 9324 11118 9336
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 11790 9324 11796 9376
rect 11848 9364 11854 9376
rect 12066 9364 12072 9376
rect 11848 9336 12072 9364
rect 11848 9324 11854 9336
rect 12066 9324 12072 9336
rect 12124 9324 12130 9376
rect 12452 9364 12480 9404
rect 12989 9401 13001 9435
rect 13035 9432 13047 9435
rect 13078 9432 13084 9444
rect 13035 9404 13084 9432
rect 13035 9401 13047 9404
rect 12989 9395 13047 9401
rect 13078 9392 13084 9404
rect 13136 9392 13142 9444
rect 12710 9364 12716 9376
rect 12452 9336 12716 9364
rect 12710 9324 12716 9336
rect 12768 9324 12774 9376
rect 12805 9367 12863 9373
rect 12805 9333 12817 9367
rect 12851 9364 12863 9367
rect 12894 9364 12900 9376
rect 12851 9336 12900 9364
rect 12851 9333 12863 9336
rect 12805 9327 12863 9333
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 13722 9324 13728 9376
rect 13780 9324 13786 9376
rect 13832 9364 13860 9472
rect 15010 9460 15016 9472
rect 15068 9460 15074 9512
rect 15672 9500 15700 9540
rect 16666 9528 16672 9580
rect 16724 9528 16730 9580
rect 17678 9528 17684 9580
rect 17736 9528 17742 9580
rect 15838 9500 15844 9512
rect 15672 9472 15844 9500
rect 15838 9460 15844 9472
rect 15896 9460 15902 9512
rect 15930 9460 15936 9512
rect 15988 9500 15994 9512
rect 16945 9503 17003 9509
rect 16945 9500 16957 9503
rect 15988 9472 16957 9500
rect 15988 9460 15994 9472
rect 16945 9469 16957 9472
rect 16991 9469 17003 9503
rect 16945 9463 17003 9469
rect 14458 9392 14464 9444
rect 14516 9432 14522 9444
rect 14645 9435 14703 9441
rect 14645 9432 14657 9435
rect 14516 9404 14657 9432
rect 14516 9392 14522 9404
rect 14645 9401 14657 9404
rect 14691 9401 14703 9435
rect 15194 9432 15200 9444
rect 14645 9395 14703 9401
rect 14752 9404 15200 9432
rect 14752 9364 14780 9404
rect 15194 9392 15200 9404
rect 15252 9392 15258 9444
rect 13832 9336 14780 9364
rect 15378 9324 15384 9376
rect 15436 9364 15442 9376
rect 16390 9364 16396 9376
rect 15436 9336 16396 9364
rect 15436 9324 15442 9336
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 17034 9324 17040 9376
rect 17092 9364 17098 9376
rect 17773 9367 17831 9373
rect 17773 9364 17785 9367
rect 17092 9336 17785 9364
rect 17092 9324 17098 9336
rect 17773 9333 17785 9336
rect 17819 9333 17831 9367
rect 17773 9327 17831 9333
rect 1104 9274 18400 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 18400 9274
rect 1104 9200 18400 9222
rect 2314 9120 2320 9172
rect 2372 9120 2378 9172
rect 2682 9120 2688 9172
rect 2740 9160 2746 9172
rect 2777 9163 2835 9169
rect 2777 9160 2789 9163
rect 2740 9132 2789 9160
rect 2740 9120 2746 9132
rect 2777 9129 2789 9132
rect 2823 9160 2835 9163
rect 2958 9160 2964 9172
rect 2823 9132 2964 9160
rect 2823 9129 2835 9132
rect 2777 9123 2835 9129
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 3259 9163 3317 9169
rect 3259 9129 3271 9163
rect 3305 9160 3317 9163
rect 3305 9132 3648 9160
rect 3305 9129 3317 9132
rect 3259 9123 3317 9129
rect 2406 9052 2412 9104
rect 2464 9092 2470 9104
rect 3421 9095 3479 9101
rect 2464 9064 3128 9092
rect 2464 9052 2470 9064
rect 3100 9024 3128 9064
rect 3421 9061 3433 9095
rect 3467 9061 3479 9095
rect 3421 9055 3479 9061
rect 3436 9024 3464 9055
rect 3100 8996 3464 9024
rect 1670 8916 1676 8968
rect 1728 8916 1734 8968
rect 1762 8916 1768 8968
rect 1820 8956 1826 8968
rect 2498 8956 2504 8968
rect 1820 8928 2504 8956
rect 1820 8916 1826 8928
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8956 2651 8959
rect 2866 8956 2872 8968
rect 2639 8928 2872 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3620 8956 3648 9132
rect 4430 9120 4436 9172
rect 4488 9160 4494 9172
rect 6181 9163 6239 9169
rect 6181 9160 6193 9163
rect 4488 9132 6193 9160
rect 4488 9120 4494 9132
rect 6181 9129 6193 9132
rect 6227 9129 6239 9163
rect 6181 9123 6239 9129
rect 7650 9120 7656 9172
rect 7708 9160 7714 9172
rect 7745 9163 7803 9169
rect 7745 9160 7757 9163
rect 7708 9132 7757 9160
rect 7708 9120 7714 9132
rect 7745 9129 7757 9132
rect 7791 9129 7803 9163
rect 7745 9123 7803 9129
rect 9490 9120 9496 9172
rect 9548 9120 9554 9172
rect 11606 9120 11612 9172
rect 11664 9160 11670 9172
rect 14369 9163 14427 9169
rect 14369 9160 14381 9163
rect 11664 9132 14381 9160
rect 11664 9120 11670 9132
rect 14369 9129 14381 9132
rect 14415 9129 14427 9163
rect 14369 9123 14427 9129
rect 14458 9120 14464 9172
rect 14516 9160 14522 9172
rect 16850 9160 16856 9172
rect 14516 9132 16856 9160
rect 14516 9120 14522 9132
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 3786 9052 3792 9104
rect 3844 9052 3850 9104
rect 3878 9052 3884 9104
rect 3936 9092 3942 9104
rect 4341 9095 4399 9101
rect 4341 9092 4353 9095
rect 3936 9064 4353 9092
rect 3936 9052 3942 9064
rect 4341 9061 4353 9064
rect 4387 9092 4399 9095
rect 5074 9092 5080 9104
rect 4387 9064 5080 9092
rect 4387 9061 4399 9064
rect 4341 9055 4399 9061
rect 5074 9052 5080 9064
rect 5132 9092 5138 9104
rect 5994 9092 6000 9104
rect 5132 9064 6000 9092
rect 5132 9052 5138 9064
rect 5994 9052 6000 9064
rect 6052 9052 6058 9104
rect 7098 9052 7104 9104
rect 7156 9092 7162 9104
rect 8018 9092 8024 9104
rect 7156 9064 8024 9092
rect 7156 9052 7162 9064
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 9030 9052 9036 9104
rect 9088 9092 9094 9104
rect 11790 9092 11796 9104
rect 9088 9064 11796 9092
rect 9088 9052 9094 9064
rect 11790 9052 11796 9064
rect 11848 9052 11854 9104
rect 12710 9052 12716 9104
rect 12768 9092 12774 9104
rect 13630 9092 13636 9104
rect 12768 9064 13636 9092
rect 12768 9052 12774 9064
rect 13630 9052 13636 9064
rect 13688 9052 13694 9104
rect 13998 9052 14004 9104
rect 14056 9092 14062 9104
rect 15013 9095 15071 9101
rect 15013 9092 15025 9095
rect 14056 9064 15025 9092
rect 14056 9052 14062 9064
rect 15013 9061 15025 9064
rect 15059 9061 15071 9095
rect 15013 9055 15071 9061
rect 15286 9052 15292 9104
rect 15344 9092 15350 9104
rect 15930 9092 15936 9104
rect 15344 9064 15936 9092
rect 15344 9052 15350 9064
rect 15930 9052 15936 9064
rect 15988 9052 15994 9104
rect 6365 9027 6423 9033
rect 6365 9024 6377 9027
rect 4080 8996 6377 9024
rect 4080 8968 4108 8996
rect 6365 8993 6377 8996
rect 6411 8993 6423 9027
rect 7466 9024 7472 9036
rect 6365 8987 6423 8993
rect 6840 8996 7472 9024
rect 3786 8956 3792 8968
rect 3620 8928 3792 8956
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 4062 8916 4068 8968
rect 4120 8916 4126 8968
rect 4154 8916 4160 8968
rect 4212 8916 4218 8968
rect 4246 8916 4252 8968
rect 4304 8916 4310 8968
rect 4525 8959 4583 8965
rect 4525 8925 4537 8959
rect 4571 8956 4583 8959
rect 4890 8956 4896 8968
rect 4571 8928 4896 8956
rect 4571 8925 4583 8928
rect 4525 8919 4583 8925
rect 4890 8916 4896 8928
rect 4948 8916 4954 8968
rect 6181 8959 6239 8965
rect 6181 8925 6193 8959
rect 6227 8925 6239 8959
rect 6181 8919 6239 8925
rect 2774 8848 2780 8900
rect 2832 8848 2838 8900
rect 3050 8848 3056 8900
rect 3108 8848 3114 8900
rect 4985 8891 5043 8897
rect 4985 8857 4997 8891
rect 5031 8888 5043 8891
rect 5534 8888 5540 8900
rect 5031 8860 5540 8888
rect 5031 8857 5043 8860
rect 4985 8851 5043 8857
rect 5534 8848 5540 8860
rect 5592 8848 5598 8900
rect 6196 8888 6224 8919
rect 6454 8916 6460 8968
rect 6512 8916 6518 8968
rect 6546 8916 6552 8968
rect 6604 8916 6610 8968
rect 6840 8888 6868 8996
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 9674 9024 9680 9036
rect 9232 8996 9680 9024
rect 6914 8916 6920 8968
rect 6972 8956 6978 8968
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 6972 8928 7573 8956
rect 6972 8916 6978 8928
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 8110 8916 8116 8968
rect 8168 8916 8174 8968
rect 9232 8965 9260 8996
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 10870 9024 10876 9036
rect 9784 8996 10876 9024
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 9306 8916 9312 8968
rect 9364 8956 9370 8968
rect 9784 8965 9812 8996
rect 10870 8984 10876 8996
rect 10928 9024 10934 9036
rect 13648 9024 13676 9052
rect 14274 9024 14280 9036
rect 10928 8996 12204 9024
rect 13648 8996 14280 9024
rect 10928 8984 10934 8996
rect 9585 8959 9643 8965
rect 9585 8956 9597 8959
rect 9364 8928 9597 8956
rect 9364 8916 9370 8928
rect 9585 8925 9597 8928
rect 9631 8925 9643 8959
rect 9585 8919 9643 8925
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 9858 8916 9864 8968
rect 9916 8916 9922 8968
rect 9950 8916 9956 8968
rect 10008 8956 10014 8968
rect 10045 8959 10103 8965
rect 10045 8956 10057 8959
rect 10008 8928 10057 8956
rect 10008 8916 10014 8928
rect 10045 8925 10057 8928
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8956 10195 8959
rect 10410 8956 10416 8968
rect 10183 8928 10416 8956
rect 10183 8925 10195 8928
rect 10137 8919 10195 8925
rect 6196 8860 6868 8888
rect 7006 8848 7012 8900
rect 7064 8888 7070 8900
rect 7064 8860 7880 8888
rect 7064 8848 7070 8860
rect 1026 8780 1032 8832
rect 1084 8820 1090 8832
rect 1489 8823 1547 8829
rect 1489 8820 1501 8823
rect 1084 8792 1501 8820
rect 1084 8780 1090 8792
rect 1489 8789 1501 8792
rect 1535 8789 1547 8823
rect 1489 8783 1547 8789
rect 3142 8780 3148 8832
rect 3200 8820 3206 8832
rect 3253 8823 3311 8829
rect 3253 8820 3265 8823
rect 3200 8792 3265 8820
rect 3200 8780 3206 8792
rect 3253 8789 3265 8792
rect 3299 8789 3311 8823
rect 3253 8783 3311 8789
rect 4614 8780 4620 8832
rect 4672 8820 4678 8832
rect 4798 8820 4804 8832
rect 4672 8792 4804 8820
rect 4672 8780 4678 8792
rect 4798 8780 4804 8792
rect 4856 8820 4862 8832
rect 5077 8823 5135 8829
rect 5077 8820 5089 8823
rect 4856 8792 5089 8820
rect 4856 8780 4862 8792
rect 5077 8789 5089 8792
rect 5123 8789 5135 8823
rect 5552 8820 5580 8848
rect 6822 8820 6828 8832
rect 5552 8792 6828 8820
rect 5077 8783 5135 8789
rect 6822 8780 6828 8792
rect 6880 8820 6886 8832
rect 7377 8823 7435 8829
rect 7377 8820 7389 8823
rect 6880 8792 7389 8820
rect 6880 8780 6886 8792
rect 7377 8789 7389 8792
rect 7423 8789 7435 8823
rect 7852 8820 7880 8860
rect 7926 8848 7932 8900
rect 7984 8848 7990 8900
rect 9493 8891 9551 8897
rect 9493 8857 9505 8891
rect 9539 8888 9551 8891
rect 10152 8888 10180 8919
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 11330 8956 11336 8968
rect 10744 8928 11336 8956
rect 10744 8916 10750 8928
rect 11330 8916 11336 8928
rect 11388 8956 11394 8968
rect 12176 8965 12204 8996
rect 14274 8984 14280 8996
rect 14332 8984 14338 9036
rect 14384 8996 15700 9024
rect 11793 8959 11851 8965
rect 11793 8956 11805 8959
rect 11388 8928 11805 8956
rect 11388 8916 11394 8928
rect 11793 8925 11805 8928
rect 11839 8925 11851 8959
rect 11793 8919 11851 8925
rect 12161 8959 12219 8965
rect 12161 8925 12173 8959
rect 12207 8925 12219 8959
rect 12161 8919 12219 8925
rect 9539 8860 10180 8888
rect 9539 8857 9551 8860
rect 9493 8851 9551 8857
rect 11698 8848 11704 8900
rect 11756 8888 11762 8900
rect 11885 8891 11943 8897
rect 11885 8888 11897 8891
rect 11756 8860 11897 8888
rect 11756 8848 11762 8860
rect 11885 8857 11897 8860
rect 11931 8857 11943 8891
rect 11885 8851 11943 8857
rect 11977 8891 12035 8897
rect 11977 8857 11989 8891
rect 12023 8857 12035 8891
rect 12176 8888 12204 8919
rect 12250 8916 12256 8968
rect 12308 8916 12314 8968
rect 14384 8888 14412 8996
rect 15672 8968 15700 8996
rect 14458 8916 14464 8968
rect 14516 8916 14522 8968
rect 14734 8916 14740 8968
rect 14792 8916 14798 8968
rect 14829 8959 14887 8965
rect 14829 8925 14841 8959
rect 14875 8956 14887 8959
rect 14918 8956 14924 8968
rect 14875 8928 14924 8956
rect 14875 8925 14887 8928
rect 14829 8919 14887 8925
rect 14918 8916 14924 8928
rect 14976 8916 14982 8968
rect 15197 8959 15255 8965
rect 15197 8925 15209 8959
rect 15243 8956 15255 8959
rect 15243 8928 15516 8956
rect 15243 8925 15255 8928
rect 15197 8919 15255 8925
rect 12176 8860 14412 8888
rect 11977 8851 12035 8857
rect 8662 8820 8668 8832
rect 7852 8792 8668 8820
rect 7377 8783 7435 8789
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 9309 8823 9367 8829
rect 9309 8789 9321 8823
rect 9355 8820 9367 8823
rect 9582 8820 9588 8832
rect 9355 8792 9588 8820
rect 9355 8789 9367 8792
rect 9309 8783 9367 8789
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 11146 8780 11152 8832
rect 11204 8820 11210 8832
rect 11609 8823 11667 8829
rect 11609 8820 11621 8823
rect 11204 8792 11621 8820
rect 11204 8780 11210 8792
rect 11609 8789 11621 8792
rect 11655 8789 11667 8823
rect 11992 8820 12020 8851
rect 12526 8820 12532 8832
rect 11992 8792 12532 8820
rect 11609 8783 11667 8789
rect 12526 8780 12532 8792
rect 12584 8820 12590 8832
rect 13078 8820 13084 8832
rect 12584 8792 13084 8820
rect 12584 8780 12590 8792
rect 13078 8780 13084 8792
rect 13136 8780 13142 8832
rect 14182 8780 14188 8832
rect 14240 8780 14246 8832
rect 14366 8780 14372 8832
rect 14424 8820 14430 8832
rect 15381 8823 15439 8829
rect 15381 8820 15393 8823
rect 14424 8792 15393 8820
rect 14424 8780 14430 8792
rect 15381 8789 15393 8792
rect 15427 8789 15439 8823
rect 15488 8820 15516 8928
rect 15654 8916 15660 8968
rect 15712 8916 15718 8968
rect 15841 8959 15899 8965
rect 15841 8925 15853 8959
rect 15887 8956 15899 8959
rect 15948 8956 15976 9052
rect 15887 8928 15976 8956
rect 15887 8925 15899 8928
rect 15841 8919 15899 8925
rect 16114 8916 16120 8968
rect 16172 8916 16178 8968
rect 16206 8916 16212 8968
rect 16264 8956 16270 8968
rect 16301 8959 16359 8965
rect 16301 8956 16313 8959
rect 16264 8928 16313 8956
rect 16264 8916 16270 8928
rect 16301 8925 16313 8928
rect 16347 8925 16359 8959
rect 16301 8919 16359 8925
rect 16390 8916 16396 8968
rect 16448 8956 16454 8968
rect 16577 8959 16635 8965
rect 16577 8956 16589 8959
rect 16448 8928 16589 8956
rect 16448 8916 16454 8928
rect 16577 8925 16589 8928
rect 16623 8925 16635 8959
rect 16577 8919 16635 8925
rect 17034 8916 17040 8968
rect 17092 8916 17098 8968
rect 17402 8916 17408 8968
rect 17460 8916 17466 8968
rect 15672 8888 15700 8916
rect 15672 8860 16712 8888
rect 15654 8820 15660 8832
rect 15488 8792 15660 8820
rect 15381 8783 15439 8789
rect 15654 8780 15660 8792
rect 15712 8780 15718 8832
rect 15930 8780 15936 8832
rect 15988 8780 15994 8832
rect 16684 8829 16712 8860
rect 16669 8823 16727 8829
rect 16669 8789 16681 8823
rect 16715 8789 16727 8823
rect 16669 8783 16727 8789
rect 1104 8730 18400 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 18400 8730
rect 1104 8656 18400 8678
rect 4062 8576 4068 8628
rect 4120 8576 4126 8628
rect 4246 8576 4252 8628
rect 4304 8616 4310 8628
rect 6365 8619 6423 8625
rect 4304 8588 6316 8616
rect 4304 8576 4310 8588
rect 5718 8548 5724 8560
rect 4356 8520 5724 8548
rect 4356 8489 4384 8520
rect 5718 8508 5724 8520
rect 5776 8508 5782 8560
rect 5810 8508 5816 8560
rect 5868 8508 5874 8560
rect 5994 8508 6000 8560
rect 6052 8508 6058 8560
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 4614 8480 4620 8492
rect 4479 8452 4620 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 5166 8440 5172 8492
rect 5224 8480 5230 8492
rect 5353 8483 5411 8489
rect 5353 8480 5365 8483
rect 5224 8452 5365 8480
rect 5224 8440 5230 8452
rect 5353 8449 5365 8452
rect 5399 8449 5411 8483
rect 5537 8483 5595 8489
rect 5537 8480 5549 8483
rect 5353 8443 5411 8449
rect 5460 8452 5549 8480
rect 5460 8344 5488 8452
rect 5537 8449 5549 8452
rect 5583 8449 5595 8483
rect 5537 8443 5595 8449
rect 5721 8415 5779 8421
rect 5721 8381 5733 8415
rect 5767 8412 5779 8415
rect 5902 8412 5908 8424
rect 5767 8384 5908 8412
rect 5767 8381 5779 8384
rect 5721 8375 5779 8381
rect 5902 8372 5908 8384
rect 5960 8412 5966 8424
rect 6086 8412 6092 8424
rect 5960 8384 6092 8412
rect 5960 8372 5966 8384
rect 6086 8372 6092 8384
rect 6144 8372 6150 8424
rect 3988 8316 5488 8344
rect 3988 8288 4016 8316
rect 6178 8304 6184 8356
rect 6236 8304 6242 8356
rect 3970 8236 3976 8288
rect 4028 8236 4034 8288
rect 4433 8279 4491 8285
rect 4433 8245 4445 8279
rect 4479 8276 4491 8279
rect 4798 8276 4804 8288
rect 4479 8248 4804 8276
rect 4479 8245 4491 8248
rect 4433 8239 4491 8245
rect 4798 8236 4804 8248
rect 4856 8236 4862 8288
rect 6288 8276 6316 8588
rect 6365 8585 6377 8619
rect 6411 8616 6423 8619
rect 6411 8588 10088 8616
rect 6411 8585 6423 8588
rect 6365 8579 6423 8585
rect 6914 8508 6920 8560
rect 6972 8548 6978 8560
rect 6972 8520 7420 8548
rect 6972 8508 6978 8520
rect 6546 8440 6552 8492
rect 6604 8440 6610 8492
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8480 6791 8483
rect 7006 8480 7012 8492
rect 6779 8452 7012 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 7392 8489 7420 8520
rect 7484 8520 7788 8548
rect 7376 8483 7434 8489
rect 7376 8449 7388 8483
rect 7422 8449 7434 8483
rect 7376 8443 7434 8449
rect 6638 8372 6644 8424
rect 6696 8372 6702 8424
rect 6825 8415 6883 8421
rect 6825 8381 6837 8415
rect 6871 8412 6883 8415
rect 7098 8412 7104 8424
rect 6871 8384 7104 8412
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 7193 8415 7251 8421
rect 7193 8381 7205 8415
rect 7239 8381 7251 8415
rect 7193 8375 7251 8381
rect 7208 8344 7236 8375
rect 7282 8372 7288 8424
rect 7340 8372 7346 8424
rect 7484 8412 7512 8520
rect 7760 8492 7788 8520
rect 8478 8508 8484 8560
rect 8536 8548 8542 8560
rect 9950 8548 9956 8560
rect 8536 8520 9352 8548
rect 8536 8508 8542 8520
rect 7650 8440 7656 8492
rect 7708 8440 7714 8492
rect 7742 8440 7748 8492
rect 7800 8480 7806 8492
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 7800 8452 7849 8480
rect 7800 8440 7806 8452
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 7926 8440 7932 8492
rect 7984 8480 7990 8492
rect 8113 8483 8171 8489
rect 8113 8480 8125 8483
rect 7984 8452 8125 8480
rect 7984 8440 7990 8452
rect 8113 8449 8125 8452
rect 8159 8480 8171 8483
rect 8159 8452 8340 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 8312 8412 8340 8452
rect 8386 8440 8392 8492
rect 8444 8440 8450 8492
rect 8570 8440 8576 8492
rect 8628 8440 8634 8492
rect 8662 8440 8668 8492
rect 8720 8440 8726 8492
rect 8846 8440 8852 8492
rect 8904 8440 8910 8492
rect 9030 8440 9036 8492
rect 9088 8440 9094 8492
rect 9214 8440 9220 8492
rect 9272 8440 9278 8492
rect 9324 8489 9352 8520
rect 9416 8520 9956 8548
rect 9416 8489 9444 8520
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 10060 8548 10088 8588
rect 11330 8576 11336 8628
rect 11388 8616 11394 8628
rect 13262 8616 13268 8628
rect 11388 8588 13268 8616
rect 11388 8576 11394 8588
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 13630 8576 13636 8628
rect 13688 8616 13694 8628
rect 13688 8588 14412 8616
rect 13688 8576 13694 8588
rect 14384 8560 14412 8588
rect 14458 8576 14464 8628
rect 14516 8576 14522 8628
rect 14734 8576 14740 8628
rect 14792 8616 14798 8628
rect 14921 8619 14979 8625
rect 14921 8616 14933 8619
rect 14792 8588 14933 8616
rect 14792 8576 14798 8588
rect 14921 8585 14933 8588
rect 14967 8585 14979 8619
rect 15470 8616 15476 8628
rect 14921 8579 14979 8585
rect 15028 8588 15476 8616
rect 11517 8551 11575 8557
rect 11517 8548 11529 8551
rect 10060 8520 10180 8548
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8449 9367 8483
rect 9309 8443 9367 8449
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 9490 8440 9496 8492
rect 9548 8480 9554 8492
rect 10152 8489 10180 8520
rect 10888 8520 11529 8548
rect 10045 8483 10103 8489
rect 10045 8480 10057 8483
rect 9548 8452 10057 8480
rect 9548 8440 9554 8452
rect 10045 8449 10057 8452
rect 10091 8449 10103 8483
rect 10045 8443 10103 8449
rect 10137 8483 10195 8489
rect 10137 8449 10149 8483
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 10226 8440 10232 8492
rect 10284 8440 10290 8492
rect 10410 8440 10416 8492
rect 10468 8440 10474 8492
rect 10686 8440 10692 8492
rect 10744 8480 10750 8492
rect 10888 8489 10916 8520
rect 11517 8517 11529 8520
rect 11563 8517 11575 8551
rect 12250 8548 12256 8560
rect 11517 8511 11575 8517
rect 11808 8520 12256 8548
rect 10781 8483 10839 8489
rect 10781 8480 10793 8483
rect 10744 8452 10793 8480
rect 10744 8440 10750 8452
rect 10781 8449 10793 8452
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8449 10931 8483
rect 10873 8443 10931 8449
rect 11054 8440 11060 8492
rect 11112 8440 11118 8492
rect 11146 8440 11152 8492
rect 11204 8440 11210 8492
rect 11330 8440 11336 8492
rect 11388 8440 11394 8492
rect 11808 8489 11836 8520
rect 12250 8508 12256 8520
rect 12308 8508 12314 8560
rect 12802 8508 12808 8560
rect 12860 8508 12866 8560
rect 13173 8551 13231 8557
rect 13173 8517 13185 8551
rect 13219 8548 13231 8551
rect 13219 8520 14320 8548
rect 13219 8517 13231 8520
rect 13173 8511 13231 8517
rect 11773 8483 11836 8489
rect 11773 8480 11785 8483
rect 11762 8449 11785 8480
rect 11819 8452 11836 8483
rect 11819 8449 11831 8452
rect 11762 8443 11831 8449
rect 11762 8412 11790 8443
rect 11882 8440 11888 8492
rect 11940 8440 11946 8492
rect 11998 8483 12056 8489
rect 11998 8449 12010 8483
rect 12044 8449 12056 8483
rect 11998 8446 12056 8449
rect 12161 8483 12219 8489
rect 12161 8449 12173 8483
rect 12207 8480 12219 8483
rect 12434 8480 12440 8492
rect 12207 8452 12440 8480
rect 12207 8449 12219 8452
rect 11998 8443 12112 8446
rect 12161 8443 12219 8449
rect 12008 8418 12112 8443
rect 12434 8440 12440 8452
rect 12492 8480 12498 8492
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12492 8452 13001 8480
rect 12492 8440 12498 8452
rect 12989 8449 13001 8452
rect 13035 8480 13047 8483
rect 13449 8483 13507 8489
rect 13449 8480 13461 8483
rect 13035 8452 13461 8480
rect 13035 8449 13047 8452
rect 12989 8443 13047 8449
rect 13449 8449 13461 8452
rect 13495 8480 13507 8483
rect 13630 8480 13636 8492
rect 13495 8452 13636 8480
rect 13495 8449 13507 8452
rect 13449 8443 13507 8449
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 14292 8489 14320 8520
rect 14366 8508 14372 8560
rect 14424 8548 14430 8560
rect 15028 8548 15056 8588
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 16114 8576 16120 8628
rect 16172 8616 16178 8628
rect 16669 8619 16727 8625
rect 16669 8616 16681 8619
rect 16172 8588 16681 8616
rect 16172 8576 16178 8588
rect 16669 8585 16681 8588
rect 16715 8585 16727 8619
rect 16669 8579 16727 8585
rect 15930 8548 15936 8560
rect 14424 8520 15056 8548
rect 15120 8520 15936 8548
rect 14424 8508 14430 8520
rect 14752 8489 14780 8520
rect 14185 8483 14243 8489
rect 14185 8480 14197 8483
rect 13780 8452 14197 8480
rect 13780 8440 13786 8452
rect 14185 8449 14197 8452
rect 14231 8449 14243 8483
rect 14185 8443 14243 8449
rect 14277 8483 14335 8489
rect 14277 8449 14289 8483
rect 14323 8449 14335 8483
rect 14277 8443 14335 8449
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8449 14611 8483
rect 14553 8443 14611 8449
rect 14737 8483 14795 8489
rect 14737 8449 14749 8483
rect 14783 8449 14795 8483
rect 14737 8443 14795 8449
rect 7391 8384 7512 8412
rect 7668 8384 8248 8412
rect 8312 8384 11790 8412
rect 7391 8344 7419 8384
rect 7208 8316 7419 8344
rect 7466 8304 7472 8356
rect 7524 8344 7530 8356
rect 7561 8347 7619 8353
rect 7561 8344 7573 8347
rect 7524 8316 7573 8344
rect 7524 8304 7530 8316
rect 7561 8313 7573 8316
rect 7607 8313 7619 8347
rect 7561 8307 7619 8313
rect 7668 8276 7696 8384
rect 7745 8347 7803 8353
rect 7745 8313 7757 8347
rect 7791 8344 7803 8347
rect 7929 8347 7987 8353
rect 7791 8316 7880 8344
rect 7791 8313 7803 8316
rect 7745 8307 7803 8313
rect 6288 8248 7696 8276
rect 7852 8276 7880 8316
rect 7929 8313 7941 8347
rect 7975 8344 7987 8347
rect 8018 8344 8024 8356
rect 7975 8316 8024 8344
rect 7975 8313 7987 8316
rect 7929 8307 7987 8313
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 8220 8353 8248 8384
rect 8205 8347 8263 8353
rect 8205 8313 8217 8347
rect 8251 8313 8263 8347
rect 8205 8307 8263 8313
rect 8297 8347 8355 8353
rect 8297 8313 8309 8347
rect 8343 8344 8355 8347
rect 8757 8347 8815 8353
rect 8757 8344 8769 8347
rect 8343 8316 8769 8344
rect 8343 8313 8355 8316
rect 8297 8307 8355 8313
rect 8757 8313 8769 8316
rect 8803 8313 8815 8347
rect 9582 8344 9588 8356
rect 8757 8307 8815 8313
rect 8864 8316 9588 8344
rect 8110 8276 8116 8288
rect 7852 8248 8116 8276
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 8220 8276 8248 8307
rect 8864 8276 8892 8316
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 9674 8304 9680 8356
rect 9732 8304 9738 8356
rect 9766 8304 9772 8356
rect 9824 8304 9830 8356
rect 10502 8304 10508 8356
rect 10560 8344 10566 8356
rect 12084 8344 12112 8418
rect 13262 8372 13268 8424
rect 13320 8412 13326 8424
rect 13541 8415 13599 8421
rect 13541 8412 13553 8415
rect 13320 8384 13553 8412
rect 13320 8372 13326 8384
rect 13541 8381 13553 8384
rect 13587 8381 13599 8415
rect 13541 8375 13599 8381
rect 13998 8372 14004 8424
rect 14056 8372 14062 8424
rect 14093 8415 14151 8421
rect 14093 8381 14105 8415
rect 14139 8412 14151 8415
rect 14366 8412 14372 8424
rect 14139 8384 14372 8412
rect 14139 8381 14151 8384
rect 14093 8375 14151 8381
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 14568 8412 14596 8443
rect 14826 8440 14832 8492
rect 14884 8440 14890 8492
rect 15120 8489 15148 8520
rect 15930 8508 15936 8520
rect 15988 8508 15994 8560
rect 16574 8548 16580 8560
rect 16316 8520 16580 8548
rect 15105 8483 15163 8489
rect 15105 8449 15117 8483
rect 15151 8449 15163 8483
rect 15105 8443 15163 8449
rect 15194 8440 15200 8492
rect 15252 8440 15258 8492
rect 15286 8440 15292 8492
rect 15344 8440 15350 8492
rect 15473 8483 15531 8489
rect 15473 8449 15485 8483
rect 15519 8449 15531 8483
rect 15473 8443 15531 8449
rect 15565 8483 15623 8489
rect 15565 8449 15577 8483
rect 15611 8480 15623 8483
rect 15746 8480 15752 8492
rect 15611 8452 15752 8480
rect 15611 8449 15623 8452
rect 15565 8443 15623 8449
rect 15488 8412 15516 8443
rect 15746 8440 15752 8452
rect 15804 8440 15810 8492
rect 15838 8440 15844 8492
rect 15896 8440 15902 8492
rect 16114 8440 16120 8492
rect 16172 8440 16178 8492
rect 16316 8489 16344 8520
rect 16574 8508 16580 8520
rect 16632 8508 16638 8560
rect 17034 8548 17040 8560
rect 16868 8520 17040 8548
rect 16301 8483 16359 8489
rect 16301 8449 16313 8483
rect 16347 8449 16359 8483
rect 16301 8443 16359 8449
rect 16482 8440 16488 8492
rect 16540 8440 16546 8492
rect 16868 8489 16896 8520
rect 17034 8508 17040 8520
rect 17092 8508 17098 8560
rect 16853 8483 16911 8489
rect 16853 8449 16865 8483
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 16942 8440 16948 8492
rect 17000 8440 17006 8492
rect 15657 8415 15715 8421
rect 15657 8412 15669 8415
rect 14568 8384 15669 8412
rect 15657 8381 15669 8384
rect 15703 8381 15715 8415
rect 15657 8375 15715 8381
rect 16025 8415 16083 8421
rect 16025 8381 16037 8415
rect 16071 8412 16083 8415
rect 16393 8415 16451 8421
rect 16393 8412 16405 8415
rect 16071 8384 16405 8412
rect 16071 8381 16083 8384
rect 16025 8375 16083 8381
rect 16393 8381 16405 8384
rect 16439 8381 16451 8415
rect 16393 8375 16451 8381
rect 10560 8316 12112 8344
rect 10560 8304 10566 8316
rect 13354 8304 13360 8356
rect 13412 8344 13418 8356
rect 13633 8347 13691 8353
rect 13633 8344 13645 8347
rect 13412 8316 13645 8344
rect 13412 8304 13418 8316
rect 13633 8313 13645 8316
rect 13679 8313 13691 8347
rect 13633 8307 13691 8313
rect 14642 8304 14648 8356
rect 14700 8344 14706 8356
rect 15933 8347 15991 8353
rect 15933 8344 15945 8347
rect 14700 8316 15945 8344
rect 14700 8304 14706 8316
rect 15933 8313 15945 8316
rect 15979 8313 15991 8347
rect 15933 8307 15991 8313
rect 8220 8248 8892 8276
rect 9490 8236 9496 8288
rect 9548 8276 9554 8288
rect 10686 8276 10692 8288
rect 9548 8248 10692 8276
rect 9548 8236 9554 8248
rect 10686 8236 10692 8248
rect 10744 8276 10750 8288
rect 12158 8276 12164 8288
rect 10744 8248 12164 8276
rect 10744 8236 10750 8248
rect 12158 8236 12164 8248
rect 12216 8276 12222 8288
rect 12618 8276 12624 8288
rect 12216 8248 12624 8276
rect 12216 8236 12222 8248
rect 12618 8236 12624 8248
rect 12676 8236 12682 8288
rect 13265 8279 13323 8285
rect 13265 8245 13277 8279
rect 13311 8276 13323 8279
rect 13722 8276 13728 8288
rect 13311 8248 13728 8276
rect 13311 8245 13323 8248
rect 13265 8239 13323 8245
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 13906 8236 13912 8288
rect 13964 8276 13970 8288
rect 14553 8279 14611 8285
rect 14553 8276 14565 8279
rect 13964 8248 14565 8276
rect 13964 8236 13970 8248
rect 14553 8245 14565 8248
rect 14599 8245 14611 8279
rect 14553 8239 14611 8245
rect 14734 8236 14740 8288
rect 14792 8276 14798 8288
rect 15746 8276 15752 8288
rect 14792 8248 15752 8276
rect 14792 8236 14798 8248
rect 15746 8236 15752 8248
rect 15804 8236 15810 8288
rect 1104 8186 18400 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 18400 8186
rect 1104 8112 18400 8134
rect 2961 8075 3019 8081
rect 2961 8041 2973 8075
rect 3007 8072 3019 8075
rect 3602 8072 3608 8084
rect 3007 8044 3608 8072
rect 3007 8041 3019 8044
rect 2961 8035 3019 8041
rect 3602 8032 3608 8044
rect 3660 8032 3666 8084
rect 6457 8075 6515 8081
rect 6457 8041 6469 8075
rect 6503 8072 6515 8075
rect 6546 8072 6552 8084
rect 6503 8044 6552 8072
rect 6503 8041 6515 8044
rect 6457 8035 6515 8041
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 6822 8032 6828 8084
rect 6880 8072 6886 8084
rect 6880 8044 7328 8072
rect 6880 8032 6886 8044
rect 2869 8007 2927 8013
rect 2869 7973 2881 8007
rect 2915 8004 2927 8007
rect 4338 8004 4344 8016
rect 2915 7976 4344 8004
rect 2915 7973 2927 7976
rect 2869 7967 2927 7973
rect 4338 7964 4344 7976
rect 4396 7964 4402 8016
rect 4525 8007 4583 8013
rect 4525 7973 4537 8007
rect 4571 7973 4583 8007
rect 4525 7967 4583 7973
rect 3510 7896 3516 7948
rect 3568 7936 3574 7948
rect 4249 7939 4307 7945
rect 4249 7936 4261 7939
rect 3568 7908 4261 7936
rect 3568 7896 3574 7908
rect 4249 7905 4261 7908
rect 4295 7905 4307 7939
rect 4540 7936 4568 7967
rect 5626 7964 5632 8016
rect 5684 8004 5690 8016
rect 6086 8004 6092 8016
rect 5684 7976 6092 8004
rect 5684 7964 5690 7976
rect 6086 7964 6092 7976
rect 6144 8004 6150 8016
rect 6144 7976 6960 8004
rect 6144 7964 6150 7976
rect 5077 7939 5135 7945
rect 5077 7936 5089 7939
rect 4540 7908 5089 7936
rect 4249 7899 4307 7905
rect 5077 7905 5089 7908
rect 5123 7936 5135 7939
rect 6638 7936 6644 7948
rect 5123 7908 6644 7936
rect 5123 7905 5135 7908
rect 5077 7899 5135 7905
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 6932 7945 6960 7976
rect 6917 7939 6975 7945
rect 6917 7905 6929 7939
rect 6963 7905 6975 7939
rect 7300 7936 7328 8044
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 7469 8075 7527 8081
rect 7469 8072 7481 8075
rect 7432 8044 7481 8072
rect 7432 8032 7438 8044
rect 7469 8041 7481 8044
rect 7515 8072 7527 8075
rect 8202 8072 8208 8084
rect 7515 8044 8208 8072
rect 7515 8041 7527 8044
rect 7469 8035 7527 8041
rect 8202 8032 8208 8044
rect 8260 8072 8266 8084
rect 10502 8072 10508 8084
rect 8260 8044 10508 8072
rect 8260 8032 8266 8044
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 10594 8032 10600 8084
rect 10652 8072 10658 8084
rect 13357 8075 13415 8081
rect 10652 8044 13308 8072
rect 10652 8032 10658 8044
rect 7558 7964 7564 8016
rect 7616 8004 7622 8016
rect 9490 8004 9496 8016
rect 7616 7976 9496 8004
rect 7616 7964 7622 7976
rect 9490 7964 9496 7976
rect 9548 7964 9554 8016
rect 9582 7964 9588 8016
rect 9640 8004 9646 8016
rect 11514 8004 11520 8016
rect 9640 7976 11520 8004
rect 9640 7964 9646 7976
rect 11514 7964 11520 7976
rect 11572 7964 11578 8016
rect 12066 8004 12072 8016
rect 11808 7976 12072 8004
rect 9125 7939 9183 7945
rect 7300 7908 7420 7936
rect 6917 7899 6975 7905
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 3326 7868 3332 7880
rect 2823 7840 3332 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 3326 7828 3332 7840
rect 3384 7828 3390 7880
rect 3418 7828 3424 7880
rect 3476 7868 3482 7880
rect 3789 7871 3847 7877
rect 3789 7868 3801 7871
rect 3476 7840 3801 7868
rect 3476 7828 3482 7840
rect 3789 7837 3801 7840
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 3970 7828 3976 7880
rect 4028 7828 4034 7880
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7868 4491 7871
rect 4522 7868 4528 7880
rect 4479 7840 4528 7868
rect 4479 7837 4491 7840
rect 4433 7831 4491 7837
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 4614 7828 4620 7880
rect 4672 7868 4678 7880
rect 4798 7868 4804 7880
rect 4672 7840 4804 7868
rect 4672 7828 4678 7840
rect 3050 7760 3056 7812
rect 3108 7800 3114 7812
rect 4724 7800 4752 7840
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 5442 7828 5448 7880
rect 5500 7828 5506 7880
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 3108 7772 4752 7800
rect 3108 7760 3114 7772
rect 4065 7735 4123 7741
rect 4065 7701 4077 7735
rect 4111 7732 4123 7735
rect 4522 7732 4528 7744
rect 4111 7704 4528 7732
rect 4111 7701 4123 7704
rect 4065 7695 4123 7701
rect 4522 7692 4528 7704
rect 4580 7692 4586 7744
rect 5552 7732 5580 7831
rect 5810 7828 5816 7880
rect 5868 7828 5874 7880
rect 5994 7877 6000 7880
rect 5961 7871 6000 7877
rect 5961 7837 5973 7871
rect 5961 7831 6000 7837
rect 5994 7828 6000 7831
rect 6052 7828 6058 7880
rect 6270 7828 6276 7880
rect 6328 7877 6334 7880
rect 6328 7831 6336 7877
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7868 6791 7871
rect 6779 7840 6960 7868
rect 6779 7837 6791 7840
rect 6733 7831 6791 7837
rect 6328 7828 6334 7831
rect 5721 7803 5779 7809
rect 5721 7769 5733 7803
rect 5767 7800 5779 7803
rect 6089 7803 6147 7809
rect 6089 7800 6101 7803
rect 5767 7772 6101 7800
rect 5767 7769 5779 7772
rect 5721 7763 5779 7769
rect 6089 7769 6101 7772
rect 6135 7769 6147 7803
rect 6089 7763 6147 7769
rect 6181 7803 6239 7809
rect 6181 7769 6193 7803
rect 6227 7769 6239 7803
rect 6181 7763 6239 7769
rect 5902 7732 5908 7744
rect 5552 7704 5908 7732
rect 5902 7692 5908 7704
rect 5960 7692 5966 7744
rect 5994 7692 6000 7744
rect 6052 7732 6058 7744
rect 6196 7732 6224 7763
rect 6932 7744 6960 7840
rect 7282 7828 7288 7880
rect 7340 7828 7346 7880
rect 7392 7877 7420 7908
rect 9125 7905 9137 7939
rect 9171 7936 9183 7939
rect 9674 7936 9680 7948
rect 9171 7908 9680 7936
rect 9171 7905 9183 7908
rect 9125 7899 9183 7905
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 10502 7936 10508 7948
rect 9784 7908 10508 7936
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7837 7435 7871
rect 7377 7831 7435 7837
rect 7561 7871 7619 7877
rect 7561 7837 7573 7871
rect 7607 7868 7619 7871
rect 7834 7868 7840 7880
rect 7607 7840 7840 7868
rect 7607 7837 7619 7840
rect 7561 7831 7619 7837
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 9214 7868 9220 7880
rect 8352 7840 9220 7868
rect 8352 7828 8358 7840
rect 9214 7828 9220 7840
rect 9272 7828 9278 7880
rect 9306 7828 9312 7880
rect 9364 7828 9370 7880
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 9784 7868 9812 7908
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 11149 7939 11207 7945
rect 11149 7905 11161 7939
rect 11195 7936 11207 7939
rect 11609 7939 11667 7945
rect 11609 7936 11621 7939
rect 11195 7908 11621 7936
rect 11195 7905 11207 7908
rect 11149 7899 11207 7905
rect 11609 7905 11621 7908
rect 11655 7905 11667 7939
rect 11609 7899 11667 7905
rect 9858 7877 9864 7880
rect 9447 7840 9812 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9856 7831 9864 7877
rect 9858 7828 9864 7831
rect 9916 7828 9922 7880
rect 10042 7828 10048 7880
rect 10100 7828 10106 7880
rect 10226 7877 10232 7880
rect 10173 7871 10232 7877
rect 10173 7868 10185 7871
rect 10152 7837 10185 7868
rect 10219 7837 10232 7871
rect 10152 7831 10232 7837
rect 7300 7772 9904 7800
rect 7300 7744 7328 7772
rect 6052 7704 6224 7732
rect 6052 7692 6058 7704
rect 6362 7692 6368 7744
rect 6420 7732 6426 7744
rect 6549 7735 6607 7741
rect 6549 7732 6561 7735
rect 6420 7704 6561 7732
rect 6420 7692 6426 7704
rect 6549 7701 6561 7704
rect 6595 7701 6607 7735
rect 6549 7695 6607 7701
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7101 7735 7159 7741
rect 7101 7732 7113 7735
rect 6972 7704 7113 7732
rect 6972 7692 6978 7704
rect 7101 7701 7113 7704
rect 7147 7701 7159 7735
rect 7101 7695 7159 7701
rect 7282 7692 7288 7744
rect 7340 7692 7346 7744
rect 9490 7692 9496 7744
rect 9548 7732 9554 7744
rect 9585 7735 9643 7741
rect 9585 7732 9597 7735
rect 9548 7704 9597 7732
rect 9548 7692 9554 7704
rect 9585 7701 9597 7704
rect 9631 7701 9643 7735
rect 9585 7695 9643 7701
rect 9674 7692 9680 7744
rect 9732 7692 9738 7744
rect 9876 7732 9904 7772
rect 9950 7760 9956 7812
rect 10008 7760 10014 7812
rect 10152 7732 10180 7831
rect 10226 7828 10232 7831
rect 10284 7828 10290 7880
rect 10318 7828 10324 7880
rect 10376 7828 10382 7880
rect 11049 7871 11107 7877
rect 11049 7868 11061 7871
rect 10980 7840 11061 7868
rect 10980 7800 11008 7840
rect 11049 7837 11061 7840
rect 11095 7837 11107 7871
rect 11049 7831 11107 7837
rect 11238 7828 11244 7880
rect 11296 7828 11302 7880
rect 11330 7828 11336 7880
rect 11388 7828 11394 7880
rect 11514 7828 11520 7880
rect 11572 7828 11578 7880
rect 11808 7877 11836 7976
rect 12066 7964 12072 7976
rect 12124 7964 12130 8016
rect 12434 7964 12440 8016
rect 12492 8004 12498 8016
rect 13170 8004 13176 8016
rect 12492 7976 13176 8004
rect 12492 7964 12498 7976
rect 13170 7964 13176 7976
rect 13228 7964 13234 8016
rect 13280 8004 13308 8044
rect 13357 8041 13369 8075
rect 13403 8072 13415 8075
rect 13722 8072 13728 8084
rect 13403 8044 13728 8072
rect 13403 8041 13415 8044
rect 13357 8035 13415 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 14182 8032 14188 8084
rect 14240 8032 14246 8084
rect 15654 8032 15660 8084
rect 15712 8072 15718 8084
rect 15933 8075 15991 8081
rect 15933 8072 15945 8075
rect 15712 8044 15945 8072
rect 15712 8032 15718 8044
rect 15933 8041 15945 8044
rect 15979 8072 15991 8075
rect 16114 8072 16120 8084
rect 15979 8044 16120 8072
rect 15979 8041 15991 8044
rect 15933 8035 15991 8041
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 15286 8004 15292 8016
rect 13280 7976 15292 8004
rect 15286 7964 15292 7976
rect 15344 8004 15350 8016
rect 15746 8004 15752 8016
rect 15344 7976 15752 8004
rect 15344 7964 15350 7976
rect 15746 7964 15752 7976
rect 15804 7964 15810 8016
rect 11885 7939 11943 7945
rect 11885 7905 11897 7939
rect 11931 7936 11943 7939
rect 12158 7936 12164 7948
rect 11931 7908 12164 7936
rect 11931 7905 11943 7908
rect 11885 7899 11943 7905
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 13265 7939 13323 7945
rect 13265 7905 13277 7939
rect 13311 7936 13323 7939
rect 13630 7936 13636 7948
rect 13311 7908 13636 7936
rect 13311 7905 13323 7908
rect 13265 7899 13323 7905
rect 11793 7871 11851 7877
rect 11793 7837 11805 7871
rect 11839 7837 11851 7871
rect 11793 7831 11851 7837
rect 11974 7828 11980 7880
rect 12032 7828 12038 7880
rect 12069 7871 12127 7877
rect 12069 7837 12081 7871
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 12084 7800 12112 7831
rect 12250 7828 12256 7880
rect 12308 7828 12314 7880
rect 12618 7828 12624 7880
rect 12676 7868 12682 7880
rect 13280 7868 13308 7899
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 13725 7939 13783 7945
rect 13725 7905 13737 7939
rect 13771 7936 13783 7939
rect 13771 7908 14228 7936
rect 13771 7905 13783 7908
rect 13725 7899 13783 7905
rect 12676 7840 13308 7868
rect 12676 7828 12682 7840
rect 13538 7828 13544 7880
rect 13596 7828 13602 7880
rect 14090 7828 14096 7880
rect 14148 7828 14154 7880
rect 14200 7868 14228 7908
rect 14556 7871 14614 7877
rect 14556 7868 14568 7871
rect 14200 7840 14568 7868
rect 14556 7837 14568 7840
rect 14602 7837 14614 7871
rect 14556 7831 14614 7837
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 15749 7871 15807 7877
rect 15749 7868 15761 7871
rect 15528 7840 15761 7868
rect 15528 7828 15534 7840
rect 15749 7837 15761 7840
rect 15795 7837 15807 7871
rect 15749 7831 15807 7837
rect 15933 7871 15991 7877
rect 15933 7837 15945 7871
rect 15979 7868 15991 7871
rect 16206 7868 16212 7880
rect 15979 7840 16212 7868
rect 15979 7837 15991 7840
rect 15933 7831 15991 7837
rect 16206 7828 16212 7840
rect 16264 7828 16270 7880
rect 17773 7871 17831 7877
rect 17773 7837 17785 7871
rect 17819 7837 17831 7871
rect 17773 7831 17831 7837
rect 14642 7800 14648 7812
rect 10980 7772 11100 7800
rect 12084 7772 14648 7800
rect 9876 7704 10180 7732
rect 10873 7735 10931 7741
rect 10873 7701 10885 7735
rect 10919 7732 10931 7735
rect 10962 7732 10968 7744
rect 10919 7704 10968 7732
rect 10919 7701 10931 7704
rect 10873 7695 10931 7701
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 11072 7732 11100 7772
rect 14642 7760 14648 7772
rect 14700 7760 14706 7812
rect 17788 7800 17816 7831
rect 14752 7772 17816 7800
rect 12710 7732 12716 7744
rect 11072 7704 12716 7732
rect 12710 7692 12716 7704
rect 12768 7692 12774 7744
rect 13170 7692 13176 7744
rect 13228 7732 13234 7744
rect 14752 7741 14780 7772
rect 14553 7735 14611 7741
rect 14553 7732 14565 7735
rect 13228 7704 14565 7732
rect 13228 7692 13234 7704
rect 14553 7701 14565 7704
rect 14599 7701 14611 7735
rect 14553 7695 14611 7701
rect 14737 7735 14795 7741
rect 14737 7701 14749 7735
rect 14783 7701 14795 7735
rect 14737 7695 14795 7701
rect 15286 7692 15292 7744
rect 15344 7732 15350 7744
rect 15838 7732 15844 7744
rect 15344 7704 15844 7732
rect 15344 7692 15350 7704
rect 15838 7692 15844 7704
rect 15896 7692 15902 7744
rect 17954 7692 17960 7744
rect 18012 7692 18018 7744
rect 1104 7642 18400 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 18400 7642
rect 1104 7568 18400 7590
rect 3053 7531 3111 7537
rect 3053 7497 3065 7531
rect 3099 7528 3111 7531
rect 3234 7528 3240 7540
rect 3099 7500 3240 7528
rect 3099 7497 3111 7500
rect 3053 7491 3111 7497
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 5813 7531 5871 7537
rect 3988 7500 5764 7528
rect 2869 7463 2927 7469
rect 2869 7429 2881 7463
rect 2915 7460 2927 7463
rect 2915 7432 3556 7460
rect 2915 7429 2927 7432
rect 2869 7423 2927 7429
rect 3528 7404 3556 7432
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 3418 7392 3424 7404
rect 2547 7364 3424 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 3510 7352 3516 7404
rect 3568 7352 3574 7404
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7392 3847 7395
rect 3878 7392 3884 7404
rect 3835 7364 3884 7392
rect 3835 7361 3847 7364
rect 3789 7355 3847 7361
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 3988 7401 4016 7500
rect 5350 7460 5356 7472
rect 4356 7432 5356 7460
rect 3973 7395 4031 7401
rect 3973 7361 3985 7395
rect 4019 7361 4031 7395
rect 3973 7355 4031 7361
rect 4062 7352 4068 7404
rect 4120 7392 4126 7404
rect 4356 7401 4384 7432
rect 5350 7420 5356 7432
rect 5408 7420 5414 7472
rect 4249 7395 4307 7401
rect 4249 7392 4261 7395
rect 4120 7364 4261 7392
rect 4120 7352 4126 7364
rect 4249 7361 4261 7364
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 3234 7284 3240 7336
rect 3292 7324 3298 7336
rect 4540 7324 4568 7355
rect 4706 7352 4712 7404
rect 4764 7392 4770 7404
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 4764 7364 5641 7392
rect 4764 7352 4770 7364
rect 5629 7361 5641 7364
rect 5675 7361 5687 7395
rect 5736 7392 5764 7500
rect 5813 7497 5825 7531
rect 5859 7528 5871 7531
rect 6270 7528 6276 7540
rect 5859 7500 6276 7528
rect 5859 7497 5871 7500
rect 5813 7491 5871 7497
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 6546 7488 6552 7540
rect 6604 7528 6610 7540
rect 6914 7528 6920 7540
rect 6604 7500 6920 7528
rect 6604 7488 6610 7500
rect 6914 7488 6920 7500
rect 6972 7488 6978 7540
rect 7374 7488 7380 7540
rect 7432 7488 7438 7540
rect 7834 7488 7840 7540
rect 7892 7528 7898 7540
rect 9674 7528 9680 7540
rect 7892 7500 9680 7528
rect 7892 7488 7898 7500
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 9858 7488 9864 7540
rect 9916 7528 9922 7540
rect 10045 7531 10103 7537
rect 10045 7528 10057 7531
rect 9916 7500 10057 7528
rect 9916 7488 9922 7500
rect 10045 7497 10057 7500
rect 10091 7497 10103 7531
rect 10045 7491 10103 7497
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 11977 7531 12035 7537
rect 11977 7528 11989 7531
rect 11296 7500 11989 7528
rect 11296 7488 11302 7500
rect 11977 7497 11989 7500
rect 12023 7497 12035 7531
rect 11977 7491 12035 7497
rect 12250 7488 12256 7540
rect 12308 7528 12314 7540
rect 12308 7500 12940 7528
rect 12308 7488 12314 7500
rect 5994 7420 6000 7472
rect 6052 7460 6058 7472
rect 7282 7460 7288 7472
rect 6052 7432 7288 7460
rect 6052 7420 6058 7432
rect 7282 7420 7288 7432
rect 7340 7420 7346 7472
rect 7392 7460 7420 7488
rect 9582 7460 9588 7472
rect 7392 7432 9588 7460
rect 6546 7392 6552 7404
rect 5736 7364 6552 7392
rect 5629 7355 5687 7361
rect 3292 7296 4568 7324
rect 3292 7284 3298 7296
rect 5350 7284 5356 7336
rect 5408 7284 5414 7336
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7293 5503 7327
rect 5445 7287 5503 7293
rect 3142 7216 3148 7268
rect 3200 7256 3206 7268
rect 3510 7256 3516 7268
rect 3200 7228 3516 7256
rect 3200 7216 3206 7228
rect 3510 7216 3516 7228
rect 3568 7256 3574 7268
rect 5460 7256 5488 7287
rect 5534 7284 5540 7336
rect 5592 7284 5598 7336
rect 3568 7228 5488 7256
rect 5644 7256 5672 7355
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 7006 7352 7012 7404
rect 7064 7392 7070 7404
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 7064 7364 7389 7392
rect 7064 7352 7070 7364
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 7650 7352 7656 7404
rect 7708 7352 7714 7404
rect 7742 7352 7748 7404
rect 7800 7352 7806 7404
rect 9232 7401 9260 7432
rect 9582 7420 9588 7432
rect 9640 7420 9646 7472
rect 10873 7463 10931 7469
rect 10873 7460 10885 7463
rect 9692 7432 10885 7460
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 9490 7352 9496 7404
rect 9548 7352 9554 7404
rect 9692 7401 9720 7432
rect 10873 7429 10885 7432
rect 10919 7429 10931 7463
rect 11514 7460 11520 7472
rect 10873 7423 10931 7429
rect 11072 7432 11520 7460
rect 9677 7395 9735 7401
rect 9677 7361 9689 7395
rect 9723 7361 9735 7395
rect 9677 7355 9735 7361
rect 10226 7352 10232 7404
rect 10284 7352 10290 7404
rect 10318 7352 10324 7404
rect 10376 7352 10382 7404
rect 10413 7395 10471 7401
rect 10413 7361 10425 7395
rect 10459 7361 10471 7395
rect 10413 7355 10471 7361
rect 10551 7395 10609 7401
rect 10551 7361 10563 7395
rect 10597 7392 10609 7395
rect 10597 7364 10916 7392
rect 10597 7361 10609 7364
rect 10551 7355 10609 7361
rect 7469 7327 7527 7333
rect 7469 7293 7481 7327
rect 7515 7324 7527 7327
rect 7834 7324 7840 7336
rect 7515 7296 7840 7324
rect 7515 7293 7527 7296
rect 7469 7287 7527 7293
rect 7834 7284 7840 7296
rect 7892 7284 7898 7336
rect 9030 7284 9036 7336
rect 9088 7284 9094 7336
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7293 9459 7327
rect 9401 7287 9459 7293
rect 7006 7256 7012 7268
rect 5644 7228 7012 7256
rect 3568 7216 3574 7228
rect 7006 7216 7012 7228
rect 7064 7216 7070 7268
rect 7929 7259 7987 7265
rect 7929 7225 7941 7259
rect 7975 7256 7987 7259
rect 9309 7259 9367 7265
rect 9309 7256 9321 7259
rect 7975 7228 9321 7256
rect 7975 7225 7987 7228
rect 7929 7219 7987 7225
rect 9309 7225 9321 7228
rect 9355 7225 9367 7259
rect 9416 7256 9444 7287
rect 10042 7284 10048 7336
rect 10100 7324 10106 7336
rect 10428 7324 10456 7355
rect 10100 7296 10456 7324
rect 10100 7284 10106 7296
rect 10686 7284 10692 7336
rect 10744 7284 10750 7336
rect 10888 7324 10916 7364
rect 10962 7352 10968 7404
rect 11020 7352 11026 7404
rect 11072 7324 11100 7432
rect 11514 7420 11520 7432
rect 11572 7420 11578 7472
rect 12268 7460 12296 7488
rect 11624 7432 12296 7460
rect 12912 7460 12940 7500
rect 14090 7488 14096 7540
rect 14148 7488 14154 7540
rect 15102 7488 15108 7540
rect 15160 7488 15166 7540
rect 15841 7531 15899 7537
rect 15841 7528 15853 7531
rect 15580 7500 15853 7528
rect 14108 7460 14136 7488
rect 12912 7432 14136 7460
rect 11238 7352 11244 7404
rect 11296 7392 11302 7404
rect 11624 7392 11652 7432
rect 11296 7364 11652 7392
rect 11296 7352 11302 7364
rect 11790 7352 11796 7404
rect 11848 7352 11854 7404
rect 11974 7352 11980 7404
rect 12032 7392 12038 7404
rect 12250 7392 12256 7404
rect 12032 7364 12256 7392
rect 12032 7352 12038 7364
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 12434 7352 12440 7404
rect 12492 7352 12498 7404
rect 12618 7352 12624 7404
rect 12676 7352 12682 7404
rect 12912 7401 12940 7432
rect 14642 7420 14648 7472
rect 14700 7460 14706 7472
rect 15580 7460 15608 7500
rect 15841 7497 15853 7500
rect 15887 7497 15899 7531
rect 15841 7491 15899 7497
rect 14700 7432 15608 7460
rect 14700 7420 14706 7432
rect 12897 7395 12955 7401
rect 12897 7361 12909 7395
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 12986 7352 12992 7404
rect 13044 7352 13050 7404
rect 13170 7352 13176 7404
rect 13228 7392 13234 7404
rect 13357 7395 13415 7401
rect 13357 7392 13369 7395
rect 13228 7364 13369 7392
rect 13228 7352 13234 7364
rect 13357 7361 13369 7364
rect 13403 7361 13415 7395
rect 13357 7355 13415 7361
rect 13538 7352 13544 7404
rect 13596 7352 13602 7404
rect 13630 7352 13636 7404
rect 13688 7392 13694 7404
rect 13688 7364 13860 7392
rect 13688 7352 13694 7364
rect 10888 7296 11100 7324
rect 11146 7284 11152 7336
rect 11204 7324 11210 7336
rect 11517 7327 11575 7333
rect 11517 7324 11529 7327
rect 11204 7296 11529 7324
rect 11204 7284 11210 7296
rect 11517 7293 11529 7296
rect 11563 7293 11575 7327
rect 11517 7287 11575 7293
rect 12802 7284 12808 7336
rect 12860 7284 12866 7336
rect 13832 7333 13860 7364
rect 13906 7352 13912 7404
rect 13964 7352 13970 7404
rect 13998 7352 14004 7404
rect 14056 7392 14062 7404
rect 14093 7395 14151 7401
rect 14093 7392 14105 7395
rect 14056 7364 14105 7392
rect 14056 7352 14062 7364
rect 14093 7361 14105 7364
rect 14139 7392 14151 7395
rect 14182 7392 14188 7404
rect 14139 7364 14188 7392
rect 14139 7361 14151 7364
rect 14093 7355 14151 7361
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 15286 7352 15292 7404
rect 15344 7352 15350 7404
rect 15580 7401 15608 7432
rect 15565 7395 15623 7401
rect 15565 7361 15577 7395
rect 15611 7361 15623 7395
rect 15565 7355 15623 7361
rect 15746 7352 15752 7404
rect 15804 7352 15810 7404
rect 16206 7352 16212 7404
rect 16264 7352 16270 7404
rect 16942 7352 16948 7404
rect 17000 7392 17006 7404
rect 17221 7395 17279 7401
rect 17221 7392 17233 7395
rect 17000 7364 17233 7392
rect 17000 7352 17006 7364
rect 17221 7361 17233 7364
rect 17267 7361 17279 7395
rect 17221 7355 17279 7361
rect 13081 7327 13139 7333
rect 13081 7293 13093 7327
rect 13127 7293 13139 7327
rect 13081 7287 13139 7293
rect 13265 7327 13323 7333
rect 13265 7293 13277 7327
rect 13311 7324 13323 7327
rect 13725 7327 13783 7333
rect 13725 7324 13737 7327
rect 13311 7296 13737 7324
rect 13311 7293 13323 7296
rect 13265 7287 13323 7293
rect 13725 7293 13737 7296
rect 13771 7293 13783 7327
rect 13725 7287 13783 7293
rect 13817 7327 13875 7333
rect 13817 7293 13829 7327
rect 13863 7324 13875 7327
rect 14734 7324 14740 7336
rect 13863 7296 14740 7324
rect 13863 7293 13875 7296
rect 13817 7287 13875 7293
rect 12529 7259 12587 7265
rect 9416 7228 12434 7256
rect 9309 7219 9367 7225
rect 2866 7148 2872 7200
rect 2924 7148 2930 7200
rect 3329 7191 3387 7197
rect 3329 7157 3341 7191
rect 3375 7188 3387 7191
rect 3694 7188 3700 7200
rect 3375 7160 3700 7188
rect 3375 7157 3387 7160
rect 3329 7151 3387 7157
rect 3694 7148 3700 7160
rect 3752 7148 3758 7200
rect 3786 7148 3792 7200
rect 3844 7188 3850 7200
rect 4065 7191 4123 7197
rect 4065 7188 4077 7191
rect 3844 7160 4077 7188
rect 3844 7148 3850 7160
rect 4065 7157 4077 7160
rect 4111 7157 4123 7191
rect 4065 7151 4123 7157
rect 4338 7148 4344 7200
rect 4396 7188 4402 7200
rect 5626 7188 5632 7200
rect 4396 7160 5632 7188
rect 4396 7148 4402 7160
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 11146 7188 11152 7200
rect 6512 7160 11152 7188
rect 6512 7148 6518 7160
rect 11146 7148 11152 7160
rect 11204 7148 11210 7200
rect 11422 7148 11428 7200
rect 11480 7188 11486 7200
rect 11609 7191 11667 7197
rect 11609 7188 11621 7191
rect 11480 7160 11621 7188
rect 11480 7148 11486 7160
rect 11609 7157 11621 7160
rect 11655 7157 11667 7191
rect 12406 7188 12434 7228
rect 12529 7225 12541 7259
rect 12575 7256 12587 7259
rect 13096 7256 13124 7287
rect 14734 7284 14740 7296
rect 14792 7284 14798 7336
rect 15194 7284 15200 7336
rect 15252 7324 15258 7336
rect 15473 7327 15531 7333
rect 15473 7324 15485 7327
rect 15252 7296 15485 7324
rect 15252 7284 15258 7296
rect 15473 7293 15485 7296
rect 15519 7293 15531 7327
rect 15473 7287 15531 7293
rect 16117 7327 16175 7333
rect 16117 7293 16129 7327
rect 16163 7324 16175 7327
rect 16390 7324 16396 7336
rect 16163 7296 16396 7324
rect 16163 7293 16175 7296
rect 16117 7287 16175 7293
rect 12575 7228 13124 7256
rect 12575 7225 12587 7228
rect 12529 7219 12587 7225
rect 13354 7216 13360 7268
rect 13412 7256 13418 7268
rect 15381 7259 15439 7265
rect 15381 7256 15393 7259
rect 13412 7228 15393 7256
rect 13412 7216 13418 7228
rect 14366 7188 14372 7200
rect 12406 7160 14372 7188
rect 11609 7151 11667 7157
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 14734 7148 14740 7200
rect 14792 7188 14798 7200
rect 14844 7188 14872 7228
rect 15381 7225 15393 7228
rect 15427 7225 15439 7259
rect 16132 7256 16160 7287
rect 16390 7284 16396 7296
rect 16448 7284 16454 7336
rect 16850 7284 16856 7336
rect 16908 7324 16914 7336
rect 17037 7327 17095 7333
rect 17037 7324 17049 7327
rect 16908 7296 17049 7324
rect 16908 7284 16914 7296
rect 17037 7293 17049 7296
rect 17083 7293 17095 7327
rect 17037 7287 17095 7293
rect 15381 7219 15439 7225
rect 15488 7228 16160 7256
rect 14792 7160 14872 7188
rect 14792 7148 14798 7160
rect 15194 7148 15200 7200
rect 15252 7188 15258 7200
rect 15488 7188 15516 7228
rect 15252 7160 15516 7188
rect 15252 7148 15258 7160
rect 15562 7148 15568 7200
rect 15620 7188 15626 7200
rect 16025 7191 16083 7197
rect 16025 7188 16037 7191
rect 15620 7160 16037 7188
rect 15620 7148 15626 7160
rect 16025 7157 16037 7160
rect 16071 7157 16083 7191
rect 16025 7151 16083 7157
rect 1104 7098 18400 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 18400 7098
rect 1104 7024 18400 7046
rect 2866 6944 2872 6996
rect 2924 6984 2930 6996
rect 5534 6984 5540 6996
rect 2924 6956 5540 6984
rect 2924 6944 2930 6956
rect 5534 6944 5540 6956
rect 5592 6944 5598 6996
rect 7009 6987 7067 6993
rect 7009 6953 7021 6987
rect 7055 6984 7067 6987
rect 7742 6984 7748 6996
rect 7055 6956 7748 6984
rect 7055 6953 7067 6956
rect 7009 6947 7067 6953
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 9858 6944 9864 6996
rect 9916 6984 9922 6996
rect 10594 6984 10600 6996
rect 9916 6956 10600 6984
rect 9916 6944 9922 6956
rect 10594 6944 10600 6956
rect 10652 6944 10658 6996
rect 12710 6984 12716 6996
rect 11808 6956 12716 6984
rect 6273 6919 6331 6925
rect 6273 6916 6285 6919
rect 5552 6888 6285 6916
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 5552 6848 5580 6888
rect 6273 6885 6285 6888
rect 6319 6885 6331 6919
rect 6273 6879 6331 6885
rect 7098 6876 7104 6928
rect 7156 6916 7162 6928
rect 8110 6916 8116 6928
rect 7156 6888 8116 6916
rect 7156 6876 7162 6888
rect 8110 6876 8116 6888
rect 8168 6876 8174 6928
rect 9398 6876 9404 6928
rect 9456 6916 9462 6928
rect 11808 6916 11836 6956
rect 12710 6944 12716 6956
rect 12768 6984 12774 6996
rect 13630 6984 13636 6996
rect 12768 6956 13636 6984
rect 12768 6944 12774 6956
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 14274 6944 14280 6996
rect 14332 6984 14338 6996
rect 15746 6984 15752 6996
rect 14332 6956 15752 6984
rect 14332 6944 14338 6956
rect 15746 6944 15752 6956
rect 15804 6944 15810 6996
rect 9456 6888 11836 6916
rect 9456 6876 9462 6888
rect 11882 6876 11888 6928
rect 11940 6876 11946 6928
rect 15838 6916 15844 6928
rect 14476 6888 15844 6916
rect 5994 6848 6000 6860
rect 3476 6820 5580 6848
rect 3476 6808 3482 6820
rect 5552 6789 5580 6820
rect 5828 6820 6000 6848
rect 5445 6783 5503 6789
rect 5445 6749 5457 6783
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 5537 6783 5595 6789
rect 5537 6749 5549 6783
rect 5583 6749 5595 6783
rect 5537 6743 5595 6749
rect 5261 6647 5319 6653
rect 5261 6613 5273 6647
rect 5307 6644 5319 6647
rect 5350 6644 5356 6656
rect 5307 6616 5356 6644
rect 5307 6613 5319 6616
rect 5261 6607 5319 6613
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 5460 6644 5488 6743
rect 5718 6740 5724 6792
rect 5776 6740 5782 6792
rect 5828 6789 5856 6820
rect 5994 6808 6000 6820
rect 6052 6808 6058 6860
rect 6178 6808 6184 6860
rect 6236 6848 6242 6860
rect 10594 6848 10600 6860
rect 6236 6820 10600 6848
rect 6236 6808 6242 6820
rect 10594 6808 10600 6820
rect 10652 6848 10658 6860
rect 11422 6848 11428 6860
rect 10652 6820 11428 6848
rect 10652 6808 10658 6820
rect 11422 6808 11428 6820
rect 11480 6848 11486 6860
rect 11698 6848 11704 6860
rect 11480 6820 11704 6848
rect 11480 6808 11486 6820
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 11790 6808 11796 6860
rect 11848 6848 11854 6860
rect 14185 6851 14243 6857
rect 14185 6848 14197 6851
rect 11848 6820 14197 6848
rect 11848 6808 11854 6820
rect 14185 6817 14197 6820
rect 14231 6817 14243 6851
rect 14476 6848 14504 6888
rect 15838 6876 15844 6888
rect 15896 6876 15902 6928
rect 16577 6919 16635 6925
rect 16577 6885 16589 6919
rect 16623 6916 16635 6919
rect 16850 6916 16856 6928
rect 16623 6888 16856 6916
rect 16623 6885 16635 6888
rect 16577 6879 16635 6885
rect 16850 6876 16856 6888
rect 16908 6876 16914 6928
rect 14185 6811 14243 6817
rect 14384 6820 14504 6848
rect 14553 6851 14611 6857
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6780 7067 6783
rect 7098 6780 7104 6792
rect 7055 6752 7104 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 7285 6783 7343 6789
rect 7285 6749 7297 6783
rect 7331 6749 7343 6783
rect 7285 6743 7343 6749
rect 5997 6715 6055 6721
rect 5997 6681 6009 6715
rect 6043 6712 6055 6715
rect 6546 6712 6552 6724
rect 6043 6684 6552 6712
rect 6043 6681 6055 6684
rect 5997 6675 6055 6681
rect 6546 6672 6552 6684
rect 6604 6672 6610 6724
rect 7193 6715 7251 6721
rect 7193 6712 7205 6715
rect 7117 6684 7205 6712
rect 6270 6644 6276 6656
rect 5460 6616 6276 6644
rect 6270 6604 6276 6616
rect 6328 6644 6334 6656
rect 6638 6644 6644 6656
rect 6328 6616 6644 6644
rect 6328 6604 6334 6616
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 6822 6604 6828 6656
rect 6880 6644 6886 6656
rect 7117 6644 7145 6684
rect 7193 6681 7205 6684
rect 7239 6681 7251 6715
rect 7300 6712 7328 6743
rect 7374 6740 7380 6792
rect 7432 6740 7438 6792
rect 7561 6783 7619 6789
rect 7561 6749 7573 6783
rect 7607 6780 7619 6783
rect 7653 6783 7711 6789
rect 7653 6780 7665 6783
rect 7607 6752 7665 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 7653 6749 7665 6752
rect 7699 6780 7711 6783
rect 7742 6780 7748 6792
rect 7699 6752 7748 6780
rect 7699 6749 7711 6752
rect 7653 6743 7711 6749
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6780 7895 6783
rect 8202 6780 8208 6792
rect 7883 6752 8208 6780
rect 7883 6749 7895 6752
rect 7837 6743 7895 6749
rect 8202 6740 8208 6752
rect 8260 6780 8266 6792
rect 10042 6780 10048 6792
rect 8260 6752 10048 6780
rect 8260 6740 8266 6752
rect 10042 6740 10048 6752
rect 10100 6780 10106 6792
rect 10778 6780 10784 6792
rect 10100 6752 10784 6780
rect 10100 6740 10106 6752
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 11330 6740 11336 6792
rect 11388 6780 11394 6792
rect 11885 6783 11943 6789
rect 11885 6780 11897 6783
rect 11388 6752 11897 6780
rect 11388 6740 11394 6752
rect 11885 6749 11897 6752
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 11974 6740 11980 6792
rect 12032 6780 12038 6792
rect 12069 6783 12127 6789
rect 12069 6780 12081 6783
rect 12032 6752 12081 6780
rect 12032 6740 12038 6752
rect 12069 6749 12081 6752
rect 12115 6780 12127 6783
rect 13814 6780 13820 6792
rect 12115 6752 13820 6780
rect 12115 6749 12127 6752
rect 12069 6743 12127 6749
rect 13814 6740 13820 6752
rect 13872 6740 13878 6792
rect 14384 6789 14412 6820
rect 14553 6817 14565 6851
rect 14599 6848 14611 6851
rect 16206 6848 16212 6860
rect 14599 6820 16212 6848
rect 14599 6817 14611 6820
rect 14553 6811 14611 6817
rect 14369 6783 14427 6789
rect 14369 6749 14381 6783
rect 14415 6749 14427 6783
rect 14369 6743 14427 6749
rect 14458 6740 14464 6792
rect 14516 6740 14522 6792
rect 14645 6783 14703 6789
rect 14645 6749 14657 6783
rect 14691 6780 14703 6783
rect 14918 6780 14924 6792
rect 14691 6752 14924 6780
rect 14691 6749 14703 6752
rect 14645 6743 14703 6749
rect 14918 6740 14924 6752
rect 14976 6740 14982 6792
rect 15102 6740 15108 6792
rect 15160 6740 15166 6792
rect 15212 6789 15240 6820
rect 16206 6808 16212 6820
rect 16264 6848 16270 6860
rect 16393 6851 16451 6857
rect 16393 6848 16405 6851
rect 16264 6820 16405 6848
rect 16264 6808 16270 6820
rect 16393 6817 16405 6820
rect 16439 6817 16451 6851
rect 16393 6811 16451 6817
rect 15197 6783 15255 6789
rect 15197 6749 15209 6783
rect 15243 6749 15255 6783
rect 15197 6743 15255 6749
rect 15286 6740 15292 6792
rect 15344 6740 15350 6792
rect 15470 6740 15476 6792
rect 15528 6740 15534 6792
rect 7469 6715 7527 6721
rect 7469 6712 7481 6715
rect 7300 6684 7481 6712
rect 7193 6675 7251 6681
rect 7469 6681 7481 6684
rect 7515 6681 7527 6715
rect 7469 6675 7527 6681
rect 8110 6672 8116 6724
rect 8168 6712 8174 6724
rect 10962 6712 10968 6724
rect 8168 6684 10968 6712
rect 8168 6672 8174 6684
rect 10962 6672 10968 6684
rect 11020 6672 11026 6724
rect 16853 6715 16911 6721
rect 16853 6681 16865 6715
rect 16899 6712 16911 6715
rect 16942 6712 16948 6724
rect 16899 6684 16948 6712
rect 16899 6681 16911 6684
rect 16853 6675 16911 6681
rect 16942 6672 16948 6684
rect 17000 6712 17006 6724
rect 17678 6712 17684 6724
rect 17000 6684 17684 6712
rect 17000 6672 17006 6684
rect 17678 6672 17684 6684
rect 17736 6672 17742 6724
rect 6880 6616 7145 6644
rect 6880 6604 6886 6616
rect 7650 6604 7656 6656
rect 7708 6644 7714 6656
rect 7745 6647 7803 6653
rect 7745 6644 7757 6647
rect 7708 6616 7757 6644
rect 7708 6604 7714 6616
rect 7745 6613 7757 6616
rect 7791 6613 7803 6647
rect 7745 6607 7803 6613
rect 12158 6604 12164 6656
rect 12216 6644 12222 6656
rect 13538 6644 13544 6656
rect 12216 6616 13544 6644
rect 12216 6604 12222 6616
rect 13538 6604 13544 6616
rect 13596 6604 13602 6656
rect 14550 6604 14556 6656
rect 14608 6644 14614 6656
rect 14829 6647 14887 6653
rect 14829 6644 14841 6647
rect 14608 6616 14841 6644
rect 14608 6604 14614 6616
rect 14829 6613 14841 6616
rect 14875 6613 14887 6647
rect 14829 6607 14887 6613
rect 1104 6554 18400 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 18400 6554
rect 1104 6480 18400 6502
rect 6178 6440 6184 6452
rect 4908 6412 6184 6440
rect 2866 6332 2872 6384
rect 2924 6332 2930 6384
rect 3085 6375 3143 6381
rect 3085 6341 3097 6375
rect 3131 6372 3143 6375
rect 3329 6375 3387 6381
rect 3329 6372 3341 6375
rect 3131 6344 3341 6372
rect 3131 6341 3143 6344
rect 3085 6335 3143 6341
rect 3329 6341 3341 6344
rect 3375 6341 3387 6375
rect 3329 6335 3387 6341
rect 3697 6375 3755 6381
rect 3697 6341 3709 6375
rect 3743 6372 3755 6375
rect 3743 6344 4292 6372
rect 3743 6341 3755 6344
rect 3697 6335 3755 6341
rect 3510 6264 3516 6316
rect 3568 6264 3574 6316
rect 3786 6264 3792 6316
rect 3844 6264 3850 6316
rect 4264 6313 4292 6344
rect 4908 6335 4936 6412
rect 6178 6400 6184 6412
rect 6236 6400 6242 6452
rect 6822 6400 6828 6452
rect 6880 6440 6886 6452
rect 7098 6440 7104 6452
rect 6880 6412 7104 6440
rect 6880 6400 6886 6412
rect 7098 6400 7104 6412
rect 7156 6440 7162 6452
rect 7285 6443 7343 6449
rect 7285 6440 7297 6443
rect 7156 6412 7297 6440
rect 7156 6400 7162 6412
rect 7285 6409 7297 6412
rect 7331 6409 7343 6443
rect 8110 6440 8116 6452
rect 7285 6403 7343 6409
rect 7392 6412 8116 6440
rect 7392 6384 7420 6412
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 8849 6443 8907 6449
rect 8849 6409 8861 6443
rect 8895 6440 8907 6443
rect 10318 6440 10324 6452
rect 8895 6412 10324 6440
rect 8895 6409 8907 6412
rect 8849 6403 8907 6409
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 11882 6400 11888 6452
rect 11940 6400 11946 6452
rect 12158 6400 12164 6452
rect 12216 6400 12222 6452
rect 12250 6400 12256 6452
rect 12308 6440 12314 6452
rect 15654 6440 15660 6452
rect 12308 6412 15056 6440
rect 12308 6400 12314 6412
rect 4893 6329 4951 6335
rect 5258 6332 5264 6384
rect 5316 6372 5322 6384
rect 5316 6344 5488 6372
rect 5316 6332 5322 6344
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6273 4215 6307
rect 4157 6267 4215 6273
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6304 4307 6307
rect 4295 6276 4752 6304
rect 4893 6295 4905 6329
rect 4939 6295 4951 6329
rect 4893 6289 4951 6295
rect 4295 6273 4307 6276
rect 4249 6267 4307 6273
rect 3528 6168 3556 6264
rect 4062 6196 4068 6248
rect 4120 6196 4126 6248
rect 4172 6168 4200 6267
rect 4341 6239 4399 6245
rect 4341 6205 4353 6239
rect 4387 6236 4399 6239
rect 4387 6208 4660 6236
rect 4387 6205 4399 6208
rect 4341 6199 4399 6205
rect 4525 6171 4583 6177
rect 4525 6168 4537 6171
rect 3528 6140 4108 6168
rect 4172 6140 4537 6168
rect 3050 6060 3056 6112
rect 3108 6060 3114 6112
rect 3237 6103 3295 6109
rect 3237 6069 3249 6103
rect 3283 6100 3295 6103
rect 3694 6100 3700 6112
rect 3283 6072 3700 6100
rect 3283 6069 3295 6072
rect 3237 6063 3295 6069
rect 3694 6060 3700 6072
rect 3752 6060 3758 6112
rect 3878 6060 3884 6112
rect 3936 6060 3942 6112
rect 4080 6100 4108 6140
rect 4525 6137 4537 6140
rect 4571 6137 4583 6171
rect 4525 6131 4583 6137
rect 4632 6100 4660 6208
rect 4724 6168 4752 6276
rect 5166 6264 5172 6316
rect 5224 6264 5230 6316
rect 5350 6264 5356 6316
rect 5408 6264 5414 6316
rect 5460 6313 5488 6344
rect 5626 6332 5632 6384
rect 5684 6372 5690 6384
rect 5684 6344 6224 6372
rect 5684 6332 5690 6344
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 4801 6239 4859 6245
rect 4801 6205 4813 6239
rect 4847 6236 4859 6239
rect 5184 6236 5212 6264
rect 4847 6208 5212 6236
rect 4847 6205 4859 6208
rect 4801 6199 4859 6205
rect 5258 6196 5264 6248
rect 5316 6236 5322 6248
rect 5552 6236 5580 6267
rect 5994 6264 6000 6316
rect 6052 6264 6058 6316
rect 6196 6313 6224 6344
rect 6546 6332 6552 6384
rect 6604 6372 6610 6384
rect 6917 6375 6975 6381
rect 6917 6372 6929 6375
rect 6604 6344 6929 6372
rect 6604 6332 6610 6344
rect 6917 6341 6929 6344
rect 6963 6341 6975 6375
rect 6917 6335 6975 6341
rect 7006 6332 7012 6384
rect 7064 6372 7070 6384
rect 7374 6372 7380 6384
rect 7064 6344 7380 6372
rect 7064 6332 7070 6344
rect 7374 6332 7380 6344
rect 7432 6332 7438 6384
rect 7558 6332 7564 6384
rect 7616 6372 7622 6384
rect 9953 6375 10011 6381
rect 9953 6372 9965 6375
rect 7616 6344 9965 6372
rect 7616 6332 7622 6344
rect 9953 6341 9965 6344
rect 9999 6372 10011 6375
rect 11900 6372 11928 6400
rect 9999 6344 11836 6372
rect 11900 6344 12664 6372
rect 9999 6341 10011 6344
rect 9953 6335 10011 6341
rect 6181 6307 6239 6313
rect 6181 6273 6193 6307
rect 6227 6273 6239 6307
rect 6181 6267 6239 6273
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 6825 6307 6883 6313
rect 6825 6304 6837 6307
rect 6696 6276 6837 6304
rect 6696 6264 6702 6276
rect 6825 6273 6837 6276
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 7101 6307 7159 6313
rect 7101 6273 7113 6307
rect 7147 6273 7159 6307
rect 7101 6267 7159 6273
rect 5316 6208 5580 6236
rect 5316 6196 5322 6208
rect 5810 6196 5816 6248
rect 5868 6236 5874 6248
rect 6454 6236 6460 6248
rect 5868 6208 6460 6236
rect 5868 6196 5874 6208
rect 6454 6196 6460 6208
rect 6512 6196 6518 6248
rect 7116 6236 7144 6267
rect 7650 6264 7656 6316
rect 7708 6264 7714 6316
rect 7926 6264 7932 6316
rect 7984 6264 7990 6316
rect 8110 6264 8116 6316
rect 8168 6264 8174 6316
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 8297 6307 8355 6313
rect 8297 6304 8309 6307
rect 8260 6276 8309 6304
rect 8260 6264 8266 6276
rect 8297 6273 8309 6276
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 8570 6264 8576 6316
rect 8628 6264 8634 6316
rect 8754 6264 8760 6316
rect 8812 6264 8818 6316
rect 9033 6307 9091 6313
rect 9033 6273 9045 6307
rect 9079 6273 9091 6307
rect 9033 6267 9091 6273
rect 7745 6239 7803 6245
rect 7116 6208 7696 6236
rect 7668 6180 7696 6208
rect 7745 6205 7757 6239
rect 7791 6205 7803 6239
rect 7745 6199 7803 6205
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 8478 6236 8484 6248
rect 7883 6208 8484 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 7469 6171 7527 6177
rect 7469 6168 7481 6171
rect 4724 6140 7481 6168
rect 7469 6137 7481 6140
rect 7515 6137 7527 6171
rect 7469 6131 7527 6137
rect 7650 6128 7656 6180
rect 7708 6128 7714 6180
rect 7760 6168 7788 6199
rect 8478 6196 8484 6208
rect 8536 6196 8542 6248
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6236 8723 6239
rect 9048 6236 9076 6267
rect 9122 6264 9128 6316
rect 9180 6264 9186 6316
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 9232 6236 9260 6267
rect 9398 6264 9404 6316
rect 9456 6264 9462 6316
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 8711 6208 9076 6236
rect 9140 6208 9260 6236
rect 8711 6205 8723 6208
rect 8665 6199 8723 6205
rect 8110 6168 8116 6180
rect 7760 6140 8116 6168
rect 8110 6128 8116 6140
rect 8168 6168 8174 6180
rect 8205 6171 8263 6177
rect 8205 6168 8217 6171
rect 8168 6140 8217 6168
rect 8168 6128 8174 6140
rect 8205 6137 8217 6140
rect 8251 6137 8263 6171
rect 8205 6131 8263 6137
rect 8938 6128 8944 6180
rect 8996 6168 9002 6180
rect 9140 6168 9168 6208
rect 9306 6196 9312 6248
rect 9364 6236 9370 6248
rect 9508 6236 9536 6267
rect 9858 6264 9864 6316
rect 9916 6264 9922 6316
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6304 10195 6307
rect 10410 6304 10416 6316
rect 10183 6276 10416 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 9364 6208 9536 6236
rect 9364 6196 9370 6208
rect 9582 6196 9588 6248
rect 9640 6236 9646 6248
rect 10152 6236 10180 6267
rect 10410 6264 10416 6276
rect 10468 6264 10474 6316
rect 10594 6264 10600 6316
rect 10652 6264 10658 6316
rect 10778 6264 10784 6316
rect 10836 6264 10842 6316
rect 10873 6307 10931 6313
rect 10873 6273 10885 6307
rect 10919 6304 10931 6307
rect 11422 6304 11428 6316
rect 10919 6276 11428 6304
rect 10919 6273 10931 6276
rect 10873 6267 10931 6273
rect 11422 6264 11428 6276
rect 11480 6264 11486 6316
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6273 11575 6307
rect 11517 6267 11575 6273
rect 9640 6208 10180 6236
rect 10321 6239 10379 6245
rect 9640 6196 9646 6208
rect 10321 6205 10333 6239
rect 10367 6236 10379 6239
rect 11146 6236 11152 6248
rect 10367 6208 11152 6236
rect 10367 6205 10379 6208
rect 10321 6199 10379 6205
rect 11146 6196 11152 6208
rect 11204 6196 11210 6248
rect 10226 6168 10232 6180
rect 8996 6140 9168 6168
rect 9324 6140 10232 6168
rect 8996 6128 9002 6140
rect 4080 6072 4660 6100
rect 4890 6060 4896 6112
rect 4948 6060 4954 6112
rect 5810 6060 5816 6112
rect 5868 6060 5874 6112
rect 5994 6060 6000 6112
rect 6052 6100 6058 6112
rect 9122 6100 9128 6112
rect 6052 6072 9128 6100
rect 6052 6060 6058 6072
rect 9122 6060 9128 6072
rect 9180 6100 9186 6112
rect 9324 6100 9352 6140
rect 10226 6128 10232 6140
rect 10284 6168 10290 6180
rect 10689 6171 10747 6177
rect 10689 6168 10701 6171
rect 10284 6140 10701 6168
rect 10284 6128 10290 6140
rect 10689 6137 10701 6140
rect 10735 6137 10747 6171
rect 11532 6168 11560 6267
rect 11698 6264 11704 6316
rect 11756 6264 11762 6316
rect 11808 6313 11836 6344
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 11882 6264 11888 6316
rect 11940 6304 11946 6316
rect 12250 6304 12256 6316
rect 11940 6276 12256 6304
rect 11940 6264 11946 6276
rect 12250 6264 12256 6276
rect 12308 6264 12314 6316
rect 12526 6264 12532 6316
rect 12584 6264 12590 6316
rect 12636 6313 12664 6344
rect 14366 6332 14372 6384
rect 14424 6332 14430 6384
rect 14737 6375 14795 6381
rect 14737 6341 14749 6375
rect 14783 6372 14795 6375
rect 14921 6375 14979 6381
rect 14921 6372 14933 6375
rect 14783 6344 14933 6372
rect 14783 6341 14795 6344
rect 14737 6335 14795 6341
rect 14921 6341 14933 6344
rect 14967 6341 14979 6375
rect 14921 6335 14979 6341
rect 12621 6307 12679 6313
rect 12621 6273 12633 6307
rect 12667 6273 12679 6307
rect 12621 6267 12679 6273
rect 12713 6307 12771 6313
rect 12713 6273 12725 6307
rect 12759 6273 12771 6307
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12713 6267 12771 6273
rect 12820 6276 12909 6304
rect 12342 6196 12348 6248
rect 12400 6236 12406 6248
rect 12728 6236 12756 6267
rect 12400 6208 12756 6236
rect 12820 6236 12848 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 13170 6264 13176 6316
rect 13228 6264 13234 6316
rect 13265 6307 13323 6313
rect 13265 6273 13277 6307
rect 13311 6273 13323 6307
rect 13265 6267 13323 6273
rect 13280 6236 13308 6267
rect 13446 6264 13452 6316
rect 13504 6264 13510 6316
rect 13541 6307 13599 6313
rect 13541 6273 13553 6307
rect 13587 6304 13599 6307
rect 13722 6304 13728 6316
rect 13587 6276 13728 6304
rect 13587 6273 13599 6276
rect 13541 6267 13599 6273
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 14274 6264 14280 6316
rect 14332 6304 14338 6316
rect 14461 6307 14519 6313
rect 14461 6304 14473 6307
rect 14332 6276 14473 6304
rect 14332 6264 14338 6276
rect 14461 6273 14473 6276
rect 14507 6273 14519 6307
rect 14461 6267 14519 6273
rect 14550 6264 14556 6316
rect 14608 6264 14614 6316
rect 14829 6307 14887 6313
rect 14829 6273 14841 6307
rect 14875 6273 14887 6307
rect 15028 6304 15056 6412
rect 15212 6412 15660 6440
rect 15105 6307 15163 6313
rect 15105 6304 15117 6307
rect 15028 6276 15117 6304
rect 14829 6267 14887 6273
rect 15105 6273 15117 6276
rect 15151 6273 15163 6307
rect 15105 6267 15163 6273
rect 12820 6208 13308 6236
rect 14844 6236 14872 6267
rect 15212 6236 15240 6412
rect 15654 6400 15660 6412
rect 15712 6400 15718 6452
rect 15838 6400 15844 6452
rect 15896 6440 15902 6452
rect 16025 6443 16083 6449
rect 16025 6440 16037 6443
rect 15896 6412 16037 6440
rect 15896 6400 15902 6412
rect 16025 6409 16037 6412
rect 16071 6440 16083 6443
rect 16206 6440 16212 6452
rect 16071 6412 16212 6440
rect 16071 6409 16083 6412
rect 16025 6403 16083 6409
rect 16206 6400 16212 6412
rect 16264 6400 16270 6452
rect 17218 6400 17224 6452
rect 17276 6440 17282 6452
rect 17773 6443 17831 6449
rect 17773 6440 17785 6443
rect 17276 6412 17785 6440
rect 17276 6400 17282 6412
rect 17773 6409 17785 6412
rect 17819 6409 17831 6443
rect 17773 6403 17831 6409
rect 15289 6375 15347 6381
rect 15289 6341 15301 6375
rect 15335 6372 15347 6375
rect 15930 6372 15936 6384
rect 15335 6344 15936 6372
rect 15335 6341 15347 6344
rect 15289 6335 15347 6341
rect 15930 6332 15936 6344
rect 15988 6372 15994 6384
rect 17034 6372 17040 6384
rect 15988 6344 17040 6372
rect 15988 6332 15994 6344
rect 17034 6332 17040 6344
rect 17092 6332 17098 6384
rect 15381 6307 15439 6313
rect 15381 6273 15393 6307
rect 15427 6273 15439 6307
rect 15381 6267 15439 6273
rect 15286 6236 15292 6248
rect 14844 6208 15292 6236
rect 12400 6196 12406 6208
rect 12820 6168 12848 6208
rect 10689 6131 10747 6137
rect 10796 6140 12848 6168
rect 13280 6168 13308 6208
rect 15286 6196 15292 6208
rect 15344 6196 15350 6248
rect 14550 6168 14556 6180
rect 13280 6140 14556 6168
rect 9180 6072 9352 6100
rect 9180 6060 9186 6072
rect 9674 6060 9680 6112
rect 9732 6060 9738 6112
rect 10318 6060 10324 6112
rect 10376 6100 10382 6112
rect 10796 6100 10824 6140
rect 14550 6128 14556 6140
rect 14608 6168 14614 6180
rect 14918 6168 14924 6180
rect 14608 6140 14924 6168
rect 14608 6128 14614 6140
rect 14918 6128 14924 6140
rect 14976 6128 14982 6180
rect 10376 6072 10824 6100
rect 10376 6060 10382 6072
rect 10870 6060 10876 6112
rect 10928 6100 10934 6112
rect 11057 6103 11115 6109
rect 11057 6100 11069 6103
rect 10928 6072 11069 6100
rect 10928 6060 10934 6072
rect 11057 6069 11069 6072
rect 11103 6069 11115 6103
rect 11057 6063 11115 6069
rect 11146 6060 11152 6112
rect 11204 6100 11210 6112
rect 11974 6100 11980 6112
rect 11204 6072 11980 6100
rect 11204 6060 11210 6072
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 12250 6060 12256 6112
rect 12308 6060 12314 6112
rect 12986 6060 12992 6112
rect 13044 6060 13050 6112
rect 14458 6060 14464 6112
rect 14516 6100 14522 6112
rect 15396 6100 15424 6267
rect 15746 6264 15752 6316
rect 15804 6304 15810 6316
rect 15841 6307 15899 6313
rect 15841 6304 15853 6307
rect 15804 6276 15853 6304
rect 15804 6264 15810 6276
rect 15841 6273 15853 6276
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 16850 6264 16856 6316
rect 16908 6304 16914 6316
rect 16945 6307 17003 6313
rect 16945 6304 16957 6307
rect 16908 6276 16957 6304
rect 16908 6264 16914 6276
rect 16945 6273 16957 6276
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 17034 6196 17040 6248
rect 17092 6196 17098 6248
rect 14516 6072 15424 6100
rect 14516 6060 14522 6072
rect 1104 6010 18400 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 18400 6010
rect 1104 5936 18400 5958
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 3421 5899 3479 5905
rect 3421 5896 3433 5899
rect 2924 5868 3433 5896
rect 2924 5856 2930 5868
rect 3421 5865 3433 5868
rect 3467 5896 3479 5899
rect 3602 5896 3608 5908
rect 3467 5868 3608 5896
rect 3467 5865 3479 5868
rect 3421 5859 3479 5865
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 3694 5856 3700 5908
rect 3752 5896 3758 5908
rect 4341 5899 4399 5905
rect 4341 5896 4353 5899
rect 3752 5868 4353 5896
rect 3752 5856 3758 5868
rect 4341 5865 4353 5868
rect 4387 5865 4399 5899
rect 4341 5859 4399 5865
rect 4798 5856 4804 5908
rect 4856 5856 4862 5908
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 5166 5896 5172 5908
rect 4948 5868 5172 5896
rect 4948 5856 4954 5868
rect 5166 5856 5172 5868
rect 5224 5896 5230 5908
rect 5224 5868 5764 5896
rect 5224 5856 5230 5868
rect 5736 5828 5764 5868
rect 5810 5856 5816 5908
rect 5868 5896 5874 5908
rect 9306 5896 9312 5908
rect 5868 5868 8156 5896
rect 5868 5856 5874 5868
rect 7742 5828 7748 5840
rect 5736 5800 6132 5828
rect 3510 5760 3516 5772
rect 2746 5732 3516 5760
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 2746 5692 2774 5732
rect 3510 5720 3516 5732
rect 3568 5720 3574 5772
rect 4430 5760 4436 5772
rect 3712 5732 4436 5760
rect 3712 5692 3740 5732
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 5169 5763 5227 5769
rect 5169 5729 5181 5763
rect 5215 5760 5227 5763
rect 5534 5760 5540 5772
rect 5215 5732 5540 5760
rect 5215 5729 5227 5732
rect 5169 5723 5227 5729
rect 5534 5720 5540 5732
rect 5592 5720 5598 5772
rect 5813 5763 5871 5769
rect 5813 5729 5825 5763
rect 5859 5760 5871 5763
rect 5994 5760 6000 5772
rect 5859 5732 6000 5760
rect 5859 5729 5871 5732
rect 5813 5723 5871 5729
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 1719 5664 2774 5692
rect 3252 5664 3740 5692
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 2498 5584 2504 5636
rect 2556 5624 2562 5636
rect 3252 5633 3280 5664
rect 3878 5652 3884 5704
rect 3936 5701 3942 5704
rect 3936 5695 3972 5701
rect 3960 5661 3972 5695
rect 3936 5655 3972 5661
rect 3936 5652 3942 5655
rect 4982 5652 4988 5704
rect 5040 5652 5046 5704
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5692 5319 5695
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 5307 5664 5457 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 5629 5695 5687 5701
rect 5629 5661 5641 5695
rect 5675 5661 5687 5695
rect 5629 5655 5687 5661
rect 3237 5627 3295 5633
rect 3237 5624 3249 5627
rect 2556 5596 3249 5624
rect 2556 5584 2562 5596
rect 3237 5593 3249 5596
rect 3283 5593 3295 5627
rect 3237 5587 3295 5593
rect 3620 5596 4016 5624
rect 1486 5516 1492 5568
rect 1544 5516 1550 5568
rect 3050 5516 3056 5568
rect 3108 5556 3114 5568
rect 3620 5565 3648 5596
rect 3437 5559 3495 5565
rect 3437 5556 3449 5559
rect 3108 5528 3449 5556
rect 3108 5516 3114 5528
rect 3437 5525 3449 5528
rect 3483 5525 3495 5559
rect 3437 5519 3495 5525
rect 3605 5559 3663 5565
rect 3605 5525 3617 5559
rect 3651 5525 3663 5559
rect 3605 5519 3663 5525
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 3988 5565 4016 5596
rect 4614 5584 4620 5636
rect 4672 5624 4678 5636
rect 5166 5624 5172 5636
rect 4672 5596 5172 5624
rect 4672 5584 4678 5596
rect 5166 5584 5172 5596
rect 5224 5624 5230 5636
rect 5644 5624 5672 5655
rect 5718 5652 5724 5704
rect 5776 5692 5782 5704
rect 5776 5664 5856 5692
rect 5776 5652 5782 5664
rect 5224 5596 5672 5624
rect 5828 5624 5856 5664
rect 5902 5652 5908 5704
rect 5960 5652 5966 5704
rect 6104 5701 6132 5800
rect 7300 5800 7748 5828
rect 6454 5720 6460 5772
rect 6512 5760 6518 5772
rect 6822 5760 6828 5772
rect 6512 5732 6828 5760
rect 6512 5720 6518 5732
rect 6822 5720 6828 5732
rect 6880 5760 6886 5772
rect 7300 5769 7328 5800
rect 7742 5788 7748 5800
rect 7800 5788 7806 5840
rect 8128 5837 8156 5868
rect 8220 5868 9312 5896
rect 8113 5831 8171 5837
rect 8113 5797 8125 5831
rect 8159 5797 8171 5831
rect 8113 5791 8171 5797
rect 7285 5763 7343 5769
rect 6880 5732 6960 5760
rect 6880 5720 6886 5732
rect 6089 5695 6147 5701
rect 6089 5661 6101 5695
rect 6135 5692 6147 5695
rect 6638 5692 6644 5704
rect 6135 5664 6644 5692
rect 6135 5661 6147 5664
rect 6089 5655 6147 5661
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 6932 5701 6960 5732
rect 7285 5729 7297 5763
rect 7331 5729 7343 5763
rect 7285 5723 7343 5729
rect 7653 5763 7711 5769
rect 7653 5729 7665 5763
rect 7699 5760 7711 5763
rect 8021 5763 8079 5769
rect 8021 5760 8033 5763
rect 7699 5732 8033 5760
rect 7699 5729 7711 5732
rect 7653 5723 7711 5729
rect 8021 5729 8033 5732
rect 8067 5729 8079 5763
rect 8220 5760 8248 5868
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 9398 5856 9404 5908
rect 9456 5896 9462 5908
rect 9677 5899 9735 5905
rect 9677 5896 9689 5899
rect 9456 5868 9689 5896
rect 9456 5856 9462 5868
rect 9677 5865 9689 5868
rect 9723 5865 9735 5899
rect 11241 5899 11299 5905
rect 9677 5859 9735 5865
rect 10428 5868 11192 5896
rect 10428 5828 10456 5868
rect 8021 5723 8079 5729
rect 8128 5732 8248 5760
rect 8312 5800 10456 5828
rect 10505 5831 10563 5837
rect 6917 5695 6975 5701
rect 6917 5661 6929 5695
rect 6963 5661 6975 5695
rect 6917 5655 6975 5661
rect 7098 5652 7104 5704
rect 7156 5652 7162 5704
rect 7193 5695 7251 5701
rect 7193 5661 7205 5695
rect 7239 5661 7251 5695
rect 7193 5655 7251 5661
rect 7469 5695 7527 5701
rect 7469 5661 7481 5695
rect 7515 5692 7527 5695
rect 7558 5692 7564 5704
rect 7515 5664 7564 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 7208 5624 7236 5655
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5692 7987 5695
rect 8128 5692 8156 5732
rect 7975 5664 8156 5692
rect 7975 5661 7987 5664
rect 7929 5655 7987 5661
rect 8202 5652 8208 5704
rect 8260 5652 8266 5704
rect 5828 5596 7236 5624
rect 5224 5584 5230 5596
rect 3789 5559 3847 5565
rect 3789 5556 3801 5559
rect 3752 5528 3801 5556
rect 3752 5516 3758 5528
rect 3789 5525 3801 5528
rect 3835 5525 3847 5559
rect 3789 5519 3847 5525
rect 3973 5559 4031 5565
rect 3973 5525 3985 5559
rect 4019 5525 4031 5559
rect 3973 5519 4031 5525
rect 4982 5516 4988 5568
rect 5040 5556 5046 5568
rect 5350 5556 5356 5568
rect 5040 5528 5356 5556
rect 5040 5516 5046 5528
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 7208 5556 7236 5596
rect 7374 5584 7380 5636
rect 7432 5624 7438 5636
rect 7745 5627 7803 5633
rect 7745 5624 7757 5627
rect 7432 5596 7757 5624
rect 7432 5584 7438 5596
rect 7745 5593 7757 5596
rect 7791 5593 7803 5627
rect 7745 5587 7803 5593
rect 8312 5556 8340 5800
rect 10505 5797 10517 5831
rect 10551 5828 10563 5831
rect 11164 5828 11192 5868
rect 11241 5865 11253 5899
rect 11287 5896 11299 5899
rect 11606 5896 11612 5908
rect 11287 5868 11612 5896
rect 11287 5865 11299 5868
rect 11241 5859 11299 5865
rect 11606 5856 11612 5868
rect 11664 5856 11670 5908
rect 12253 5899 12311 5905
rect 12253 5865 12265 5899
rect 12299 5896 12311 5899
rect 12342 5896 12348 5908
rect 12299 5868 12348 5896
rect 12299 5865 12311 5868
rect 12253 5859 12311 5865
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 12529 5899 12587 5905
rect 12529 5865 12541 5899
rect 12575 5896 12587 5899
rect 13170 5896 13176 5908
rect 12575 5868 13176 5896
rect 12575 5865 12587 5868
rect 12529 5859 12587 5865
rect 13170 5856 13176 5868
rect 13228 5856 13234 5908
rect 13262 5856 13268 5908
rect 13320 5856 13326 5908
rect 15102 5896 15108 5908
rect 14660 5868 15108 5896
rect 11790 5828 11796 5840
rect 10551 5800 10732 5828
rect 11164 5800 11796 5828
rect 10551 5797 10563 5800
rect 10505 5791 10563 5797
rect 9674 5760 9680 5772
rect 8956 5732 9680 5760
rect 8478 5652 8484 5704
rect 8536 5692 8542 5704
rect 8956 5701 8984 5732
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 10226 5760 10232 5772
rect 9876 5732 10232 5760
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8536 5664 8953 5692
rect 8536 5652 8542 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 9030 5652 9036 5704
rect 9088 5690 9094 5704
rect 9125 5695 9183 5701
rect 9125 5690 9137 5695
rect 9088 5662 9137 5690
rect 9088 5652 9094 5662
rect 9125 5661 9137 5662
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5661 9275 5695
rect 9217 5655 9275 5661
rect 9309 5695 9367 5701
rect 9309 5661 9321 5695
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 8754 5584 8760 5636
rect 8812 5624 8818 5636
rect 9232 5624 9260 5655
rect 8812 5596 8984 5624
rect 8812 5584 8818 5596
rect 8956 5590 8984 5596
rect 9140 5596 9260 5624
rect 9140 5590 9168 5596
rect 8956 5562 9168 5590
rect 7208 5528 8340 5556
rect 9324 5556 9352 5655
rect 9490 5652 9496 5704
rect 9548 5652 9554 5704
rect 9876 5701 9904 5732
rect 10226 5720 10232 5732
rect 10284 5720 10290 5772
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5661 9919 5695
rect 9861 5655 9919 5661
rect 9954 5695 10012 5701
rect 9954 5661 9966 5695
rect 10000 5692 10012 5695
rect 10042 5692 10048 5704
rect 10000 5664 10048 5692
rect 10000 5661 10012 5664
rect 9954 5655 10012 5661
rect 9858 5556 9864 5568
rect 9324 5528 9864 5556
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 9968 5556 9996 5655
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 10134 5652 10140 5704
rect 10192 5652 10198 5704
rect 10318 5652 10324 5704
rect 10376 5701 10382 5704
rect 10376 5692 10384 5701
rect 10376 5664 10421 5692
rect 10376 5655 10384 5664
rect 10376 5652 10382 5655
rect 10594 5652 10600 5704
rect 10652 5652 10658 5704
rect 10704 5692 10732 5800
rect 11790 5788 11796 5800
rect 11848 5788 11854 5840
rect 12066 5788 12072 5840
rect 12124 5828 12130 5840
rect 13078 5828 13084 5840
rect 12124 5800 13084 5828
rect 12124 5788 12130 5800
rect 13078 5788 13084 5800
rect 13136 5828 13142 5840
rect 14660 5837 14688 5868
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 15746 5856 15752 5908
rect 15804 5896 15810 5908
rect 16945 5899 17003 5905
rect 16945 5896 16957 5899
rect 15804 5868 16957 5896
rect 15804 5856 15810 5868
rect 16945 5865 16957 5868
rect 16991 5865 17003 5899
rect 16945 5859 17003 5865
rect 14645 5831 14703 5837
rect 14645 5828 14657 5831
rect 13136 5800 14657 5828
rect 13136 5788 13142 5800
rect 14645 5797 14657 5800
rect 14691 5797 14703 5831
rect 14645 5791 14703 5797
rect 13173 5763 13231 5769
rect 11348 5732 12664 5760
rect 10781 5695 10839 5701
rect 10781 5692 10793 5695
rect 10704 5664 10793 5692
rect 10781 5661 10793 5664
rect 10827 5661 10839 5695
rect 10781 5655 10839 5661
rect 10870 5652 10876 5704
rect 10928 5652 10934 5704
rect 10965 5695 11023 5701
rect 10965 5661 10977 5695
rect 11011 5692 11023 5695
rect 11238 5692 11244 5704
rect 11011 5664 11244 5692
rect 11011 5661 11023 5664
rect 10965 5655 11023 5661
rect 11238 5652 11244 5664
rect 11296 5652 11302 5704
rect 10229 5627 10287 5633
rect 10229 5593 10241 5627
rect 10275 5624 10287 5627
rect 10686 5624 10692 5636
rect 10275 5596 10692 5624
rect 10275 5593 10287 5596
rect 10229 5587 10287 5593
rect 10686 5584 10692 5596
rect 10744 5584 10750 5636
rect 11348 5624 11376 5732
rect 11422 5652 11428 5704
rect 11480 5692 11486 5704
rect 11701 5695 11759 5701
rect 11701 5692 11713 5695
rect 11480 5664 11713 5692
rect 11480 5652 11486 5664
rect 11701 5661 11713 5664
rect 11747 5661 11759 5695
rect 11701 5655 11759 5661
rect 11790 5652 11796 5704
rect 11848 5652 11854 5704
rect 11974 5652 11980 5704
rect 12032 5652 12038 5704
rect 12069 5695 12127 5701
rect 12069 5661 12081 5695
rect 12115 5661 12127 5695
rect 12069 5655 12127 5661
rect 10796 5596 11376 5624
rect 10796 5556 10824 5596
rect 9968 5528 10824 5556
rect 11330 5516 11336 5568
rect 11388 5556 11394 5568
rect 12084 5556 12112 5655
rect 12434 5652 12440 5704
rect 12492 5652 12498 5704
rect 12636 5701 12664 5732
rect 13173 5729 13185 5763
rect 13219 5760 13231 5763
rect 13538 5760 13544 5772
rect 13219 5732 13544 5760
rect 13219 5729 13231 5732
rect 13173 5723 13231 5729
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 15933 5763 15991 5769
rect 14844 5732 15332 5760
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5661 12679 5695
rect 12621 5655 12679 5661
rect 12636 5624 12664 5655
rect 13630 5652 13636 5704
rect 13688 5692 13694 5704
rect 14844 5692 14872 5732
rect 13688 5664 13733 5692
rect 13832 5664 14872 5692
rect 13688 5652 13694 5664
rect 13832 5624 13860 5664
rect 14918 5652 14924 5704
rect 14976 5652 14982 5704
rect 15102 5652 15108 5704
rect 15160 5652 15166 5704
rect 15304 5701 15332 5732
rect 15933 5729 15945 5763
rect 15979 5729 15991 5763
rect 16114 5760 16120 5772
rect 15933 5723 15991 5729
rect 16040 5732 16120 5760
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5692 15347 5695
rect 15378 5692 15384 5704
rect 15335 5664 15384 5692
rect 15335 5661 15347 5664
rect 15289 5655 15347 5661
rect 15378 5652 15384 5664
rect 15436 5692 15442 5704
rect 15948 5692 15976 5723
rect 16040 5701 16068 5732
rect 16114 5720 16120 5732
rect 16172 5760 16178 5772
rect 16850 5760 16856 5772
rect 16172 5732 16856 5760
rect 16172 5720 16178 5732
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 15436 5664 15976 5692
rect 16025 5695 16083 5701
rect 15436 5652 15442 5664
rect 16025 5661 16037 5695
rect 16071 5661 16083 5695
rect 16025 5655 16083 5661
rect 16669 5695 16727 5701
rect 16669 5661 16681 5695
rect 16715 5692 16727 5695
rect 17402 5692 17408 5704
rect 16715 5664 17408 5692
rect 16715 5661 16727 5664
rect 16669 5655 16727 5661
rect 17402 5652 17408 5664
rect 17460 5652 17466 5704
rect 12636 5596 13860 5624
rect 14366 5584 14372 5636
rect 14424 5624 14430 5636
rect 14461 5627 14519 5633
rect 14461 5624 14473 5627
rect 14424 5596 14473 5624
rect 14424 5584 14430 5596
rect 14461 5593 14473 5596
rect 14507 5593 14519 5627
rect 14461 5587 14519 5593
rect 11388 5528 12112 5556
rect 11388 5516 11394 5528
rect 12894 5516 12900 5568
rect 12952 5556 12958 5568
rect 13630 5556 13636 5568
rect 12952 5528 13636 5556
rect 12952 5516 12958 5528
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 13814 5516 13820 5568
rect 13872 5516 13878 5568
rect 14476 5556 14504 5587
rect 15194 5584 15200 5636
rect 15252 5584 15258 5636
rect 16758 5624 16764 5636
rect 15396 5596 16764 5624
rect 15396 5556 15424 5596
rect 16758 5584 16764 5596
rect 16816 5584 16822 5636
rect 16853 5627 16911 5633
rect 16853 5593 16865 5627
rect 16899 5593 16911 5627
rect 16853 5587 16911 5593
rect 14476 5528 15424 5556
rect 15470 5516 15476 5568
rect 15528 5516 15534 5568
rect 16666 5516 16672 5568
rect 16724 5556 16730 5568
rect 16868 5556 16896 5587
rect 16724 5528 16896 5556
rect 16724 5516 16730 5528
rect 1104 5466 18400 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 18400 5466
rect 1104 5392 18400 5414
rect 3973 5355 4031 5361
rect 3973 5321 3985 5355
rect 4019 5352 4031 5355
rect 4062 5352 4068 5364
rect 4019 5324 4068 5352
rect 4019 5321 4031 5324
rect 3973 5315 4031 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 6822 5312 6828 5364
rect 6880 5352 6886 5364
rect 6880 5324 8156 5352
rect 6880 5312 6886 5324
rect 2038 5244 2044 5296
rect 2096 5284 2102 5296
rect 7558 5284 7564 5296
rect 2096 5256 6868 5284
rect 2096 5244 2102 5256
rect 3786 5176 3792 5228
rect 3844 5216 3850 5228
rect 4341 5219 4399 5225
rect 4341 5216 4353 5219
rect 3844 5188 4353 5216
rect 3844 5176 3850 5188
rect 4341 5185 4353 5188
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 6638 5176 6644 5228
rect 6696 5216 6702 5228
rect 6733 5219 6791 5225
rect 6733 5216 6745 5219
rect 6696 5188 6745 5216
rect 6696 5176 6702 5188
rect 6733 5185 6745 5188
rect 6779 5185 6791 5219
rect 6733 5179 6791 5185
rect 4249 5151 4307 5157
rect 4249 5117 4261 5151
rect 4295 5148 4307 5151
rect 4798 5148 4804 5160
rect 4295 5120 4804 5148
rect 4295 5117 4307 5120
rect 4249 5111 4307 5117
rect 4798 5108 4804 5120
rect 4856 5108 4862 5160
rect 6840 5148 6868 5256
rect 7024 5256 7564 5284
rect 6914 5176 6920 5228
rect 6972 5176 6978 5228
rect 7024 5225 7052 5256
rect 7558 5244 7564 5256
rect 7616 5244 7622 5296
rect 8128 5284 8156 5324
rect 8202 5312 8208 5364
rect 8260 5352 8266 5364
rect 8665 5355 8723 5361
rect 8665 5352 8677 5355
rect 8260 5324 8677 5352
rect 8260 5312 8266 5324
rect 8665 5321 8677 5324
rect 8711 5321 8723 5355
rect 8665 5315 8723 5321
rect 8754 5312 8760 5364
rect 8812 5352 8818 5364
rect 12161 5355 12219 5361
rect 8812 5324 11192 5352
rect 8812 5312 8818 5324
rect 8938 5284 8944 5296
rect 8128 5256 8944 5284
rect 8938 5244 8944 5256
rect 8996 5284 9002 5296
rect 11054 5284 11060 5296
rect 8996 5256 11060 5284
rect 8996 5244 9002 5256
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 7098 5176 7104 5228
rect 7156 5216 7162 5228
rect 8570 5216 8576 5228
rect 7156 5188 8576 5216
rect 7156 5176 7162 5188
rect 8570 5176 8576 5188
rect 8628 5176 8634 5228
rect 8846 5176 8852 5228
rect 8904 5176 8910 5228
rect 9140 5225 9168 5256
rect 11054 5244 11060 5256
rect 11112 5244 11118 5296
rect 11164 5284 11192 5324
rect 12161 5321 12173 5355
rect 12207 5352 12219 5355
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 12207 5324 13461 5352
rect 12207 5321 12219 5324
rect 12161 5315 12219 5321
rect 13449 5321 13461 5324
rect 13495 5321 13507 5355
rect 13449 5315 13507 5321
rect 13814 5312 13820 5364
rect 13872 5352 13878 5364
rect 13975 5355 14033 5361
rect 13975 5352 13987 5355
rect 13872 5324 13987 5352
rect 13872 5312 13878 5324
rect 13975 5321 13987 5324
rect 14021 5321 14033 5355
rect 14277 5355 14335 5361
rect 14277 5352 14289 5355
rect 13975 5315 14033 5321
rect 14108 5324 14289 5352
rect 13357 5287 13415 5293
rect 11164 5256 12204 5284
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 10321 5219 10379 5225
rect 10321 5185 10333 5219
rect 10367 5216 10379 5219
rect 10410 5216 10416 5228
rect 10367 5188 10416 5216
rect 10367 5185 10379 5188
rect 10321 5179 10379 5185
rect 10410 5176 10416 5188
rect 10468 5176 10474 5228
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 10781 5219 10839 5225
rect 10781 5216 10793 5219
rect 10744 5188 10793 5216
rect 10744 5176 10750 5188
rect 10781 5185 10793 5188
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 8662 5148 8668 5160
rect 6840 5120 8668 5148
rect 8662 5108 8668 5120
rect 8720 5108 8726 5160
rect 8754 5108 8760 5160
rect 8812 5108 8818 5160
rect 10505 5151 10563 5157
rect 10505 5148 10517 5151
rect 8864 5120 10517 5148
rect 4430 5040 4436 5092
rect 4488 5080 4494 5092
rect 4488 5052 5580 5080
rect 4488 5040 4494 5052
rect 4341 5015 4399 5021
rect 4341 4981 4353 5015
rect 4387 5012 4399 5015
rect 5442 5012 5448 5024
rect 4387 4984 5448 5012
rect 4387 4981 4399 4984
rect 4341 4975 4399 4981
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 5552 5012 5580 5052
rect 5626 5040 5632 5092
rect 5684 5080 5690 5092
rect 8864 5080 8892 5120
rect 10505 5117 10517 5120
rect 10551 5148 10563 5151
rect 11330 5148 11336 5160
rect 10551 5120 11336 5148
rect 10551 5117 10563 5120
rect 10505 5111 10563 5117
rect 11330 5108 11336 5120
rect 11388 5108 11394 5160
rect 12176 5157 12204 5256
rect 13357 5253 13369 5287
rect 13403 5284 13415 5287
rect 14108 5284 14136 5324
rect 14277 5321 14289 5324
rect 14323 5321 14335 5355
rect 14277 5315 14335 5321
rect 14550 5312 14556 5364
rect 14608 5352 14614 5364
rect 14608 5324 15608 5352
rect 14608 5312 14614 5324
rect 13403 5256 14136 5284
rect 13403 5253 13415 5256
rect 13357 5247 13415 5253
rect 14182 5244 14188 5296
rect 14240 5244 14246 5296
rect 15470 5244 15476 5296
rect 15528 5244 15534 5296
rect 12250 5176 12256 5228
rect 12308 5216 12314 5228
rect 12437 5219 12495 5225
rect 12437 5216 12449 5219
rect 12308 5188 12449 5216
rect 12308 5176 12314 5188
rect 12437 5185 12449 5188
rect 12483 5185 12495 5219
rect 12437 5179 12495 5185
rect 12161 5151 12219 5157
rect 12161 5117 12173 5151
rect 12207 5117 12219 5151
rect 12452 5148 12480 5179
rect 12526 5176 12532 5228
rect 12584 5176 12590 5228
rect 12710 5176 12716 5228
rect 12768 5176 12774 5228
rect 13078 5176 13084 5228
rect 13136 5216 13142 5228
rect 13265 5219 13323 5225
rect 13265 5216 13277 5219
rect 13136 5188 13277 5216
rect 13136 5176 13142 5188
rect 13265 5185 13277 5188
rect 13311 5185 13323 5219
rect 13265 5179 13323 5185
rect 13538 5176 13544 5228
rect 13596 5216 13602 5228
rect 13596 5188 14228 5216
rect 13596 5176 13602 5188
rect 12452 5120 12572 5148
rect 12161 5111 12219 5117
rect 5684 5052 8892 5080
rect 5684 5040 5690 5052
rect 9858 5040 9864 5092
rect 9916 5080 9922 5092
rect 10413 5083 10471 5089
rect 10413 5080 10425 5083
rect 9916 5052 10425 5080
rect 9916 5040 9922 5052
rect 10413 5049 10425 5052
rect 10459 5080 10471 5083
rect 10778 5080 10784 5092
rect 10459 5052 10784 5080
rect 10459 5049 10471 5052
rect 10413 5043 10471 5049
rect 10778 5040 10784 5052
rect 10836 5040 10842 5092
rect 7006 5012 7012 5024
rect 5552 4984 7012 5012
rect 7006 4972 7012 4984
rect 7064 5012 7070 5024
rect 7282 5012 7288 5024
rect 7064 4984 7288 5012
rect 7064 4972 7070 4984
rect 7282 4972 7288 4984
rect 7340 4972 7346 5024
rect 7374 4972 7380 5024
rect 7432 4972 7438 5024
rect 9033 5015 9091 5021
rect 9033 4981 9045 5015
rect 9079 5012 9091 5015
rect 10045 5015 10103 5021
rect 10045 5012 10057 5015
rect 9079 4984 10057 5012
rect 9079 4981 9091 4984
rect 9033 4975 9091 4981
rect 10045 4981 10057 4984
rect 10091 4981 10103 5015
rect 10045 4975 10103 4981
rect 10597 5015 10655 5021
rect 10597 4981 10609 5015
rect 10643 5012 10655 5015
rect 11238 5012 11244 5024
rect 10643 4984 11244 5012
rect 10643 4981 10655 4984
rect 10597 4975 10655 4981
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 12342 4972 12348 5024
rect 12400 5012 12406 5024
rect 12434 5012 12440 5024
rect 12400 4984 12440 5012
rect 12400 4972 12406 4984
rect 12434 4972 12440 4984
rect 12492 4972 12498 5024
rect 12544 5021 12572 5120
rect 13630 5108 13636 5160
rect 13688 5108 13694 5160
rect 13722 5108 13728 5160
rect 13780 5108 13786 5160
rect 14200 5148 14228 5188
rect 14274 5176 14280 5228
rect 14332 5176 14338 5228
rect 14461 5219 14519 5225
rect 14461 5185 14473 5219
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 15197 5219 15255 5225
rect 15197 5185 15209 5219
rect 15243 5185 15255 5219
rect 15197 5179 15255 5185
rect 14476 5148 14504 5179
rect 15212 5148 15240 5179
rect 15286 5176 15292 5228
rect 15344 5176 15350 5228
rect 15381 5219 15439 5225
rect 15381 5185 15393 5219
rect 15427 5216 15439 5219
rect 15488 5216 15516 5244
rect 15580 5225 15608 5324
rect 15746 5312 15752 5364
rect 15804 5352 15810 5364
rect 16393 5355 16451 5361
rect 15804 5324 16160 5352
rect 15804 5312 15810 5324
rect 16022 5284 16028 5296
rect 15856 5256 16028 5284
rect 15856 5225 15884 5256
rect 16022 5244 16028 5256
rect 16080 5244 16086 5296
rect 16132 5225 16160 5324
rect 16393 5321 16405 5355
rect 16439 5352 16451 5355
rect 16666 5352 16672 5364
rect 16439 5324 16672 5352
rect 16439 5321 16451 5324
rect 16393 5315 16451 5321
rect 16666 5312 16672 5324
rect 16724 5312 16730 5364
rect 15427 5188 15516 5216
rect 15565 5219 15623 5225
rect 15427 5185 15439 5188
rect 15381 5179 15439 5185
rect 15565 5185 15577 5219
rect 15611 5185 15623 5219
rect 15565 5179 15623 5185
rect 15841 5219 15899 5225
rect 15841 5185 15853 5219
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5185 15991 5219
rect 15933 5179 15991 5185
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5185 16175 5219
rect 16117 5179 16175 5185
rect 15657 5151 15715 5157
rect 15657 5148 15669 5151
rect 14200 5120 15056 5148
rect 15212 5120 15669 5148
rect 15028 5089 15056 5120
rect 15657 5117 15669 5120
rect 15703 5117 15715 5151
rect 15948 5148 15976 5179
rect 16206 5176 16212 5228
rect 16264 5176 16270 5228
rect 16485 5219 16543 5225
rect 16485 5216 16497 5219
rect 16408 5188 16497 5216
rect 16298 5148 16304 5160
rect 15948 5120 16304 5148
rect 15657 5111 15715 5117
rect 16298 5108 16304 5120
rect 16356 5108 16362 5160
rect 12897 5083 12955 5089
rect 12897 5049 12909 5083
rect 12943 5080 12955 5083
rect 15013 5083 15071 5089
rect 12943 5052 14044 5080
rect 12943 5049 12955 5052
rect 12897 5043 12955 5049
rect 12529 5015 12587 5021
rect 12529 4981 12541 5015
rect 12575 4981 12587 5015
rect 12529 4975 12587 4981
rect 12986 4972 12992 5024
rect 13044 4972 13050 5024
rect 13817 5015 13875 5021
rect 13817 4981 13829 5015
rect 13863 5012 13875 5015
rect 13906 5012 13912 5024
rect 13863 4984 13912 5012
rect 13863 4981 13875 4984
rect 13817 4975 13875 4981
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 14016 5021 14044 5052
rect 15013 5049 15025 5083
rect 15059 5049 15071 5083
rect 15013 5043 15071 5049
rect 15194 5040 15200 5092
rect 15252 5080 15258 5092
rect 16408 5080 16436 5188
rect 16485 5185 16497 5188
rect 16531 5185 16543 5219
rect 16485 5179 16543 5185
rect 15252 5052 16436 5080
rect 15252 5040 15258 5052
rect 14001 5015 14059 5021
rect 14001 4981 14013 5015
rect 14047 4981 14059 5015
rect 14001 4975 14059 4981
rect 1104 4922 18400 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 18400 4922
rect 1104 4848 18400 4870
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 5721 4811 5779 4817
rect 5721 4808 5733 4811
rect 5592 4780 5733 4808
rect 5592 4768 5598 4780
rect 5721 4777 5733 4780
rect 5767 4777 5779 4811
rect 8754 4808 8760 4820
rect 5721 4771 5779 4777
rect 5828 4780 8760 4808
rect 3329 4743 3387 4749
rect 3329 4709 3341 4743
rect 3375 4740 3387 4743
rect 3418 4740 3424 4752
rect 3375 4712 3424 4740
rect 3375 4709 3387 4712
rect 3329 4703 3387 4709
rect 3418 4700 3424 4712
rect 3476 4700 3482 4752
rect 5350 4700 5356 4752
rect 5408 4740 5414 4752
rect 5828 4740 5856 4780
rect 8754 4768 8760 4780
rect 8812 4808 8818 4820
rect 9950 4808 9956 4820
rect 8812 4780 9956 4808
rect 8812 4768 8818 4780
rect 9950 4768 9956 4780
rect 10008 4808 10014 4820
rect 10594 4808 10600 4820
rect 10008 4780 10600 4808
rect 10008 4768 10014 4780
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 11330 4768 11336 4820
rect 11388 4768 11394 4820
rect 11977 4811 12035 4817
rect 11977 4777 11989 4811
rect 12023 4777 12035 4811
rect 11977 4771 12035 4777
rect 12161 4811 12219 4817
rect 12161 4777 12173 4811
rect 12207 4808 12219 4811
rect 12342 4808 12348 4820
rect 12207 4780 12348 4808
rect 12207 4777 12219 4780
rect 12161 4771 12219 4777
rect 7190 4740 7196 4752
rect 5408 4712 5856 4740
rect 7024 4712 7196 4740
rect 5408 4700 5414 4712
rect 3436 4604 3464 4700
rect 5810 4672 5816 4684
rect 5644 4644 5816 4672
rect 4706 4604 4712 4616
rect 3436 4576 4712 4604
rect 4706 4564 4712 4576
rect 4764 4604 4770 4616
rect 5644 4613 5672 4644
rect 5810 4632 5816 4644
rect 5868 4672 5874 4684
rect 6549 4675 6607 4681
rect 6549 4672 6561 4675
rect 5868 4644 6561 4672
rect 5868 4632 5874 4644
rect 6549 4641 6561 4644
rect 6595 4641 6607 4675
rect 7024 4672 7052 4712
rect 7190 4700 7196 4712
rect 7248 4700 7254 4752
rect 11992 4740 12020 4771
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 13446 4768 13452 4820
rect 13504 4808 13510 4820
rect 13504 4780 14780 4808
rect 13504 4768 13510 4780
rect 14752 4752 14780 4780
rect 14826 4768 14832 4820
rect 14884 4808 14890 4820
rect 15746 4808 15752 4820
rect 14884 4780 15752 4808
rect 14884 4768 14890 4780
rect 15746 4768 15752 4780
rect 15804 4768 15810 4820
rect 15930 4768 15936 4820
rect 15988 4768 15994 4820
rect 13262 4740 13268 4752
rect 10520 4712 12020 4740
rect 12084 4712 13268 4740
rect 6549 4635 6607 4641
rect 6748 4644 7052 4672
rect 7101 4675 7159 4681
rect 5445 4607 5503 4613
rect 5445 4604 5457 4607
rect 4764 4576 5457 4604
rect 4764 4564 4770 4576
rect 5445 4573 5457 4576
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 5902 4564 5908 4616
rect 5960 4564 5966 4616
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4573 6055 4607
rect 5997 4567 6055 4573
rect 6457 4607 6515 4613
rect 6457 4573 6469 4607
rect 6503 4604 6515 4607
rect 6748 4604 6776 4644
rect 7101 4641 7113 4675
rect 7147 4672 7159 4675
rect 7653 4675 7711 4681
rect 7653 4672 7665 4675
rect 7147 4644 7665 4672
rect 7147 4641 7159 4644
rect 7101 4635 7159 4641
rect 7653 4641 7665 4644
rect 7699 4641 7711 4675
rect 7653 4635 7711 4641
rect 6503 4576 6776 4604
rect 6503 4573 6515 4576
rect 6457 4567 6515 4573
rect 2961 4539 3019 4545
rect 2961 4505 2973 4539
rect 3007 4536 3019 4539
rect 3142 4536 3148 4548
rect 3007 4508 3148 4536
rect 3007 4505 3019 4508
rect 2961 4499 3019 4505
rect 3142 4496 3148 4508
rect 3200 4496 3206 4548
rect 5261 4539 5319 4545
rect 5261 4505 5273 4539
rect 5307 4536 5319 4539
rect 5350 4536 5356 4548
rect 5307 4508 5356 4536
rect 5307 4505 5319 4508
rect 5261 4499 5319 4505
rect 5350 4496 5356 4508
rect 5408 4496 5414 4548
rect 5721 4539 5779 4545
rect 5721 4505 5733 4539
rect 5767 4505 5779 4539
rect 6012 4536 6040 4567
rect 6822 4564 6828 4616
rect 6880 4564 6886 4616
rect 6914 4564 6920 4616
rect 6972 4564 6978 4616
rect 7006 4564 7012 4616
rect 7064 4604 7070 4616
rect 7193 4607 7251 4613
rect 7193 4604 7205 4607
rect 7064 4576 7205 4604
rect 7064 4564 7070 4576
rect 7193 4573 7205 4576
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 7374 4564 7380 4616
rect 7432 4564 7438 4616
rect 7466 4564 7472 4616
rect 7524 4564 7530 4616
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4604 7803 4607
rect 7834 4604 7840 4616
rect 7791 4576 7840 4604
rect 7791 4573 7803 4576
rect 7745 4567 7803 4573
rect 7834 4564 7840 4576
rect 7892 4564 7898 4616
rect 10520 4536 10548 4712
rect 11422 4632 11428 4684
rect 11480 4672 11486 4684
rect 12084 4672 12112 4712
rect 13262 4700 13268 4712
rect 13320 4700 13326 4752
rect 14458 4740 14464 4752
rect 13556 4712 14464 4740
rect 13556 4672 13584 4712
rect 14458 4700 14464 4712
rect 14516 4700 14522 4752
rect 14734 4700 14740 4752
rect 14792 4740 14798 4752
rect 15197 4743 15255 4749
rect 15197 4740 15209 4743
rect 14792 4712 15209 4740
rect 14792 4700 14798 4712
rect 15197 4709 15209 4712
rect 15243 4709 15255 4743
rect 15197 4703 15255 4709
rect 15381 4743 15439 4749
rect 15381 4709 15393 4743
rect 15427 4740 15439 4743
rect 15427 4712 15516 4740
rect 15427 4709 15439 4712
rect 15381 4703 15439 4709
rect 11480 4644 12112 4672
rect 12406 4644 13584 4672
rect 11480 4632 11486 4644
rect 11514 4564 11520 4616
rect 11572 4564 11578 4616
rect 12406 4604 12434 4644
rect 13630 4632 13636 4684
rect 13688 4672 13694 4684
rect 15488 4672 15516 4712
rect 13688 4644 15516 4672
rect 13688 4632 13694 4644
rect 11716 4576 12434 4604
rect 6012 4508 11192 4536
rect 5721 4499 5779 4505
rect 3421 4471 3479 4477
rect 3421 4437 3433 4471
rect 3467 4468 3479 4471
rect 5626 4468 5632 4480
rect 3467 4440 5632 4468
rect 3467 4437 3479 4440
rect 3421 4431 3479 4437
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 5736 4468 5764 4499
rect 6638 4468 6644 4480
rect 5736 4440 6644 4468
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 6733 4471 6791 4477
rect 6733 4437 6745 4471
rect 6779 4468 6791 4471
rect 7098 4468 7104 4480
rect 6779 4440 7104 4468
rect 6779 4437 6791 4440
rect 6733 4431 6791 4437
rect 7098 4428 7104 4440
rect 7156 4428 7162 4480
rect 7193 4471 7251 4477
rect 7193 4437 7205 4471
rect 7239 4468 7251 4471
rect 7374 4468 7380 4480
rect 7239 4440 7380 4468
rect 7239 4437 7251 4440
rect 7193 4431 7251 4437
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 11164 4477 11192 4508
rect 11330 4496 11336 4548
rect 11388 4536 11394 4548
rect 11716 4536 11744 4576
rect 13262 4564 13268 4616
rect 13320 4564 13326 4616
rect 13446 4564 13452 4616
rect 13504 4564 13510 4616
rect 13814 4564 13820 4616
rect 13872 4564 13878 4616
rect 14369 4607 14427 4613
rect 14369 4573 14381 4607
rect 14415 4573 14427 4607
rect 15488 4604 15516 4644
rect 15654 4632 15660 4684
rect 15712 4672 15718 4684
rect 15948 4672 15976 4768
rect 15712 4644 15976 4672
rect 15712 4632 15718 4644
rect 16298 4604 16304 4616
rect 15488 4576 16304 4604
rect 14369 4567 14427 4573
rect 11388 4508 11744 4536
rect 11388 4496 11394 4508
rect 11790 4496 11796 4548
rect 11848 4496 11854 4548
rect 14090 4536 14096 4548
rect 13990 4508 14096 4536
rect 11149 4471 11207 4477
rect 11149 4437 11161 4471
rect 11195 4437 11207 4471
rect 11149 4431 11207 4437
rect 11974 4428 11980 4480
rect 12032 4477 12038 4480
rect 12032 4471 12051 4477
rect 12039 4437 12051 4471
rect 12032 4431 12051 4437
rect 12032 4428 12038 4431
rect 13354 4428 13360 4480
rect 13412 4428 13418 4480
rect 13633 4471 13691 4477
rect 13633 4437 13645 4471
rect 13679 4468 13691 4471
rect 13990 4468 14018 4508
rect 14090 4496 14096 4508
rect 14148 4536 14154 4548
rect 14384 4536 14412 4567
rect 16298 4564 16304 4576
rect 16356 4564 16362 4616
rect 14148 4508 14412 4536
rect 15933 4539 15991 4545
rect 14148 4496 14154 4508
rect 15933 4505 15945 4539
rect 15979 4536 15991 4539
rect 16114 4536 16120 4548
rect 15979 4508 16120 4536
rect 15979 4505 15991 4508
rect 15933 4499 15991 4505
rect 16114 4496 16120 4508
rect 16172 4496 16178 4548
rect 13679 4440 14018 4468
rect 13679 4437 13691 4440
rect 13633 4431 13691 4437
rect 14182 4428 14188 4480
rect 14240 4428 14246 4480
rect 1104 4378 18400 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 18400 4378
rect 1104 4304 18400 4326
rect 5721 4267 5779 4273
rect 5721 4233 5733 4267
rect 5767 4264 5779 4267
rect 5902 4264 5908 4276
rect 5767 4236 5908 4264
rect 5767 4233 5779 4236
rect 5721 4227 5779 4233
rect 5902 4224 5908 4236
rect 5960 4264 5966 4276
rect 6457 4267 6515 4273
rect 6457 4264 6469 4267
rect 5960 4236 6469 4264
rect 5960 4224 5966 4236
rect 6457 4233 6469 4236
rect 6503 4233 6515 4267
rect 6457 4227 6515 4233
rect 8570 4224 8576 4276
rect 8628 4224 8634 4276
rect 8941 4267 8999 4273
rect 8941 4233 8953 4267
rect 8987 4264 8999 4267
rect 10318 4264 10324 4276
rect 8987 4236 10324 4264
rect 8987 4233 8999 4236
rect 8941 4227 8999 4233
rect 10318 4224 10324 4236
rect 10376 4224 10382 4276
rect 10962 4224 10968 4276
rect 11020 4264 11026 4276
rect 11146 4264 11152 4276
rect 11020 4236 11152 4264
rect 11020 4224 11026 4236
rect 11146 4224 11152 4236
rect 11204 4224 11210 4276
rect 11790 4224 11796 4276
rect 11848 4264 11854 4276
rect 11848 4236 11928 4264
rect 11848 4224 11854 4236
rect 3786 4156 3792 4208
rect 3844 4156 3850 4208
rect 4706 4156 4712 4208
rect 4764 4156 4770 4208
rect 5626 4156 5632 4208
rect 5684 4196 5690 4208
rect 5997 4199 6055 4205
rect 5997 4196 6009 4199
rect 5684 4168 6009 4196
rect 5684 4156 5690 4168
rect 5997 4165 6009 4168
rect 6043 4165 6055 4199
rect 5997 4159 6055 4165
rect 6638 4156 6644 4208
rect 6696 4196 6702 4208
rect 6822 4196 6828 4208
rect 6696 4168 6828 4196
rect 6696 4156 6702 4168
rect 6822 4156 6828 4168
rect 6880 4196 6886 4208
rect 8478 4196 8484 4208
rect 6880 4168 8484 4196
rect 6880 4156 6886 4168
rect 8478 4156 8484 4168
rect 8536 4156 8542 4208
rect 8588 4196 8616 4224
rect 8757 4199 8815 4205
rect 8757 4196 8769 4199
rect 8588 4168 8769 4196
rect 8757 4165 8769 4168
rect 8803 4165 8815 4199
rect 8757 4159 8815 4165
rect 8956 4168 10088 4196
rect 8956 4140 8984 4168
rect 3142 4088 3148 4140
rect 3200 4088 3206 4140
rect 3418 4088 3424 4140
rect 3476 4088 3482 4140
rect 5353 4131 5411 4137
rect 5353 4128 5365 4131
rect 5184 4100 5365 4128
rect 5184 4069 5212 4100
rect 5353 4097 5365 4100
rect 5399 4128 5411 4131
rect 5718 4128 5724 4140
rect 5399 4100 5724 4128
rect 5399 4097 5411 4100
rect 5353 4091 5411 4097
rect 5718 4088 5724 4100
rect 5776 4088 5782 4140
rect 5810 4088 5816 4140
rect 5868 4088 5874 4140
rect 6181 4131 6239 4137
rect 6181 4097 6193 4131
rect 6227 4128 6239 4131
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 6227 4100 6377 4128
rect 6227 4097 6239 4100
rect 6181 4091 6239 4097
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 6917 4131 6975 4137
rect 6917 4097 6929 4131
rect 6963 4128 6975 4131
rect 7006 4128 7012 4140
rect 6963 4100 7012 4128
rect 6963 4097 6975 4100
rect 6917 4091 6975 4097
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 7193 4131 7251 4137
rect 7193 4097 7205 4131
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 5169 4063 5227 4069
rect 5169 4029 5181 4063
rect 5215 4029 5227 4063
rect 5169 4023 5227 4029
rect 5258 4020 5264 4072
rect 5316 4060 5322 4072
rect 5445 4063 5503 4069
rect 5445 4060 5457 4063
rect 5316 4032 5457 4060
rect 5316 4020 5322 4032
rect 5445 4029 5457 4032
rect 5491 4029 5503 4063
rect 7208 4060 7236 4091
rect 7374 4088 7380 4140
rect 7432 4088 7438 4140
rect 7745 4131 7803 4137
rect 7745 4097 7757 4131
rect 7791 4128 7803 4131
rect 8205 4131 8263 4137
rect 8205 4128 8217 4131
rect 7791 4100 8217 4128
rect 7791 4097 7803 4100
rect 7745 4091 7803 4097
rect 8205 4097 8217 4100
rect 8251 4097 8263 4131
rect 8205 4091 8263 4097
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 7561 4063 7619 4069
rect 7561 4060 7573 4063
rect 7208 4032 7573 4060
rect 5445 4023 5503 4029
rect 7561 4029 7573 4032
rect 7607 4029 7619 4063
rect 7561 4023 7619 4029
rect 7834 4020 7840 4072
rect 7892 4020 7898 4072
rect 7929 4063 7987 4069
rect 7929 4029 7941 4063
rect 7975 4029 7987 4063
rect 7929 4023 7987 4029
rect 5077 3995 5135 4001
rect 5077 3961 5089 3995
rect 5123 3992 5135 3995
rect 6641 3995 6699 4001
rect 5123 3964 5488 3992
rect 5123 3961 5135 3964
rect 5077 3955 5135 3961
rect 5460 3936 5488 3964
rect 6641 3961 6653 3995
rect 6687 3992 6699 3995
rect 6914 3992 6920 4004
rect 6687 3964 6920 3992
rect 6687 3961 6699 3964
rect 6641 3955 6699 3961
rect 6914 3952 6920 3964
rect 6972 3952 6978 4004
rect 5442 3884 5448 3936
rect 5500 3884 5506 3936
rect 5537 3927 5595 3933
rect 5537 3893 5549 3927
rect 5583 3924 5595 3927
rect 6270 3924 6276 3936
rect 5583 3896 6276 3924
rect 5583 3893 5595 3896
rect 5537 3887 5595 3893
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 6733 3927 6791 3933
rect 6733 3893 6745 3927
rect 6779 3924 6791 3927
rect 6822 3924 6828 3936
rect 6779 3896 6828 3924
rect 6779 3893 6791 3896
rect 6733 3887 6791 3893
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 7944 3924 7972 4023
rect 8018 4020 8024 4072
rect 8076 4020 8082 4072
rect 8110 4020 8116 4072
rect 8168 4060 8174 4072
rect 8680 4060 8708 4091
rect 8938 4088 8944 4140
rect 8996 4088 9002 4140
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 9125 4131 9183 4137
rect 9125 4097 9137 4131
rect 9171 4097 9183 4131
rect 9125 4091 9183 4097
rect 9048 4060 9076 4091
rect 8168 4032 9076 4060
rect 8168 4020 8174 4032
rect 9030 3952 9036 4004
rect 9088 3992 9094 4004
rect 9140 3992 9168 4091
rect 9214 4088 9220 4140
rect 9272 4088 9278 4140
rect 9324 4137 9352 4168
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 9582 4088 9588 4140
rect 9640 4088 9646 4140
rect 9766 4088 9772 4140
rect 9824 4088 9830 4140
rect 9858 4088 9864 4140
rect 9916 4088 9922 4140
rect 9953 4131 10011 4137
rect 9953 4097 9965 4131
rect 9999 4097 10011 4131
rect 10060 4128 10088 4168
rect 10686 4156 10692 4208
rect 10744 4196 10750 4208
rect 11900 4196 11928 4236
rect 11974 4224 11980 4276
rect 12032 4224 12038 4276
rect 13078 4224 13084 4276
rect 13136 4224 13142 4276
rect 13262 4224 13268 4276
rect 13320 4264 13326 4276
rect 16206 4264 16212 4276
rect 13320 4236 16212 4264
rect 13320 4224 13326 4236
rect 16206 4224 16212 4236
rect 16264 4224 16270 4276
rect 10744 4168 11836 4196
rect 11900 4168 12434 4196
rect 10744 4156 10750 4168
rect 10137 4131 10195 4137
rect 10137 4128 10149 4131
rect 10060 4100 10149 4128
rect 9953 4091 10011 4097
rect 10137 4097 10149 4100
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 9968 3992 9996 4091
rect 10502 4088 10508 4140
rect 10560 4128 10566 4140
rect 10597 4131 10655 4137
rect 10597 4128 10609 4131
rect 10560 4100 10609 4128
rect 10560 4088 10566 4100
rect 10597 4097 10609 4100
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 10778 4088 10784 4140
rect 10836 4088 10842 4140
rect 11057 4131 11115 4137
rect 11057 4097 11069 4131
rect 11103 4097 11115 4131
rect 11057 4091 11115 4097
rect 11072 4060 11100 4091
rect 11698 4088 11704 4140
rect 11756 4088 11762 4140
rect 11808 4128 11836 4168
rect 11885 4131 11943 4137
rect 11885 4128 11897 4131
rect 11808 4100 11897 4128
rect 11885 4097 11897 4100
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 11977 4131 12035 4137
rect 11977 4097 11989 4131
rect 12023 4128 12035 4131
rect 12066 4128 12072 4140
rect 12023 4100 12072 4128
rect 12023 4097 12035 4100
rect 11977 4091 12035 4097
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12158 4088 12164 4140
rect 12216 4088 12222 4140
rect 12406 4128 12434 4168
rect 13354 4156 13360 4208
rect 13412 4156 13418 4208
rect 15010 4156 15016 4208
rect 15068 4156 15074 4208
rect 16114 4196 16120 4208
rect 15948 4168 16120 4196
rect 12406 4100 13216 4128
rect 11793 4063 11851 4069
rect 11793 4060 11805 4063
rect 11072 4032 11805 4060
rect 11793 4029 11805 4032
rect 11839 4060 11851 4063
rect 12618 4060 12624 4072
rect 11839 4032 12624 4060
rect 11839 4029 11851 4032
rect 11793 4023 11851 4029
rect 12618 4020 12624 4032
rect 12676 4020 12682 4072
rect 13188 4060 13216 4100
rect 13262 4088 13268 4140
rect 13320 4088 13326 4140
rect 13449 4131 13507 4137
rect 13449 4097 13461 4131
rect 13495 4097 13507 4131
rect 13449 4091 13507 4097
rect 13464 4060 13492 4091
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 13633 4131 13691 4137
rect 13633 4128 13645 4131
rect 13596 4100 13645 4128
rect 13596 4088 13602 4100
rect 13633 4097 13645 4100
rect 13679 4097 13691 4131
rect 13633 4091 13691 4097
rect 13722 4088 13728 4140
rect 13780 4088 13786 4140
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 14921 4131 14979 4137
rect 14921 4128 14933 4131
rect 14424 4100 14933 4128
rect 14424 4088 14430 4100
rect 14921 4097 14933 4100
rect 14967 4128 14979 4131
rect 15194 4128 15200 4140
rect 14967 4100 15200 4128
rect 14967 4097 14979 4100
rect 14921 4091 14979 4097
rect 15194 4088 15200 4100
rect 15252 4088 15258 4140
rect 15654 4088 15660 4140
rect 15712 4088 15718 4140
rect 15948 4137 15976 4168
rect 16114 4156 16120 4168
rect 16172 4196 16178 4208
rect 16172 4168 16896 4196
rect 16172 4156 16178 4168
rect 15933 4131 15991 4137
rect 15933 4097 15945 4131
rect 15979 4097 15991 4131
rect 15933 4091 15991 4097
rect 16298 4088 16304 4140
rect 16356 4128 16362 4140
rect 16868 4137 16896 4168
rect 16761 4131 16819 4137
rect 16761 4128 16773 4131
rect 16356 4100 16773 4128
rect 16356 4088 16362 4100
rect 16761 4097 16773 4100
rect 16807 4097 16819 4131
rect 16761 4091 16819 4097
rect 16853 4131 16911 4137
rect 16853 4097 16865 4131
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4097 17095 4131
rect 17037 4091 17095 4097
rect 14182 4060 14188 4072
rect 13188 4032 14188 4060
rect 14182 4020 14188 4032
rect 14240 4020 14246 4072
rect 14274 4020 14280 4072
rect 14332 4060 14338 4072
rect 15672 4060 15700 4088
rect 17052 4060 17080 4091
rect 14332 4032 14964 4060
rect 15672 4032 17080 4060
rect 14332 4020 14338 4032
rect 9088 3964 9168 3992
rect 9232 3964 9996 3992
rect 10045 3995 10103 4001
rect 9088 3952 9094 3964
rect 8294 3924 8300 3936
rect 7944 3896 8300 3924
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 8754 3884 8760 3936
rect 8812 3884 8818 3936
rect 8846 3884 8852 3936
rect 8904 3924 8910 3936
rect 9232 3924 9260 3964
rect 10045 3961 10057 3995
rect 10091 3992 10103 3995
rect 10134 3992 10140 4004
rect 10091 3964 10140 3992
rect 10091 3961 10103 3964
rect 10045 3955 10103 3961
rect 10134 3952 10140 3964
rect 10192 3952 10198 4004
rect 10410 3952 10416 4004
rect 10468 3992 10474 4004
rect 14642 3992 14648 4004
rect 10468 3964 14648 3992
rect 10468 3952 10474 3964
rect 14642 3952 14648 3964
rect 14700 3952 14706 4004
rect 14936 3992 14964 4032
rect 14936 3964 16712 3992
rect 8904 3896 9260 3924
rect 9401 3927 9459 3933
rect 8904 3884 8910 3896
rect 9401 3893 9413 3927
rect 9447 3924 9459 3927
rect 9490 3924 9496 3936
rect 9447 3896 9496 3924
rect 9447 3893 9459 3896
rect 9401 3887 9459 3893
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 16574 3924 16580 3936
rect 11296 3896 16580 3924
rect 11296 3884 11302 3896
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 16684 3924 16712 3964
rect 16758 3952 16764 4004
rect 16816 3992 16822 4004
rect 16853 3995 16911 4001
rect 16853 3992 16865 3995
rect 16816 3964 16865 3992
rect 16816 3952 16822 3964
rect 16853 3961 16865 3964
rect 16899 3961 16911 3995
rect 16853 3955 16911 3961
rect 16942 3924 16948 3936
rect 16684 3896 16948 3924
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 1104 3834 18400 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 18400 3834
rect 1104 3760 18400 3782
rect 5629 3723 5687 3729
rect 5629 3689 5641 3723
rect 5675 3720 5687 3723
rect 5810 3720 5816 3732
rect 5675 3692 5816 3720
rect 5675 3689 5687 3692
rect 5629 3683 5687 3689
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 7742 3680 7748 3732
rect 7800 3680 7806 3732
rect 7834 3680 7840 3732
rect 7892 3720 7898 3732
rect 8481 3723 8539 3729
rect 8481 3720 8493 3723
rect 7892 3692 8493 3720
rect 7892 3680 7898 3692
rect 8481 3689 8493 3692
rect 8527 3689 8539 3723
rect 8481 3683 8539 3689
rect 8573 3723 8631 3729
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 8754 3720 8760 3732
rect 8619 3692 8760 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 8754 3680 8760 3692
rect 8812 3720 8818 3732
rect 9677 3723 9735 3729
rect 8812 3692 9628 3720
rect 8812 3680 8818 3692
rect 3142 3612 3148 3664
rect 3200 3652 3206 3664
rect 3200 3624 5396 3652
rect 3200 3612 3206 3624
rect 3053 3587 3111 3593
rect 3053 3553 3065 3587
rect 3099 3584 3111 3587
rect 4985 3587 5043 3593
rect 4985 3584 4997 3587
rect 3099 3556 4997 3584
rect 3099 3553 3111 3556
rect 3053 3547 3111 3553
rect 4985 3553 4997 3556
rect 5031 3584 5043 3587
rect 5258 3584 5264 3596
rect 5031 3556 5264 3584
rect 5031 3553 5043 3556
rect 4985 3547 5043 3553
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 5368 3528 5396 3624
rect 7098 3612 7104 3664
rect 7156 3652 7162 3664
rect 7469 3655 7527 3661
rect 7469 3652 7481 3655
rect 7156 3624 7481 3652
rect 7156 3612 7162 3624
rect 7469 3621 7481 3624
rect 7515 3652 7527 3655
rect 7760 3652 7788 3680
rect 9030 3652 9036 3664
rect 7515 3624 9036 3652
rect 7515 3621 7527 3624
rect 7469 3615 7527 3621
rect 9030 3612 9036 3624
rect 9088 3612 9094 3664
rect 9214 3612 9220 3664
rect 9272 3652 9278 3664
rect 9309 3655 9367 3661
rect 9309 3652 9321 3655
rect 9272 3624 9321 3652
rect 9272 3612 9278 3624
rect 9309 3621 9321 3624
rect 9355 3621 9367 3655
rect 9600 3652 9628 3692
rect 9677 3689 9689 3723
rect 9723 3720 9735 3723
rect 9858 3720 9864 3732
rect 9723 3692 9864 3720
rect 9723 3689 9735 3692
rect 9677 3683 9735 3689
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 10778 3680 10784 3732
rect 10836 3720 10842 3732
rect 11977 3723 12035 3729
rect 11977 3720 11989 3723
rect 10836 3692 11989 3720
rect 10836 3680 10842 3692
rect 11977 3689 11989 3692
rect 12023 3720 12035 3723
rect 12023 3692 12434 3720
rect 12023 3689 12035 3692
rect 11977 3683 12035 3689
rect 12161 3655 12219 3661
rect 12161 3652 12173 3655
rect 9600 3624 12173 3652
rect 9309 3615 9367 3621
rect 12161 3621 12173 3624
rect 12207 3621 12219 3655
rect 12161 3615 12219 3621
rect 6086 3544 6092 3596
rect 6144 3544 6150 3596
rect 8389 3587 8447 3593
rect 6196 3556 7420 3584
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 3436 3448 3464 3479
rect 3510 3476 3516 3528
rect 3568 3516 3574 3528
rect 3605 3519 3663 3525
rect 3605 3516 3617 3519
rect 3568 3488 3617 3516
rect 3568 3476 3574 3488
rect 3605 3485 3617 3488
rect 3651 3516 3663 3519
rect 4065 3519 4123 3525
rect 4065 3516 4077 3519
rect 3651 3488 4077 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 4065 3485 4077 3488
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 3970 3448 3976 3460
rect 3436 3420 3976 3448
rect 3970 3408 3976 3420
rect 4028 3448 4034 3460
rect 4356 3448 4384 3479
rect 5350 3476 5356 3528
rect 5408 3476 5414 3528
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 6196 3516 6224 3556
rect 5500 3488 6224 3516
rect 5500 3476 5506 3488
rect 6546 3476 6552 3528
rect 6604 3476 6610 3528
rect 6730 3476 6736 3528
rect 6788 3516 6794 3528
rect 7392 3525 7420 3556
rect 8389 3553 8401 3587
rect 8435 3584 8447 3587
rect 8478 3584 8484 3596
rect 8435 3556 8484 3584
rect 8435 3553 8447 3556
rect 8389 3547 8447 3553
rect 8478 3544 8484 3556
rect 8536 3544 8542 3596
rect 9401 3587 9459 3593
rect 9401 3584 9413 3587
rect 8680 3556 9413 3584
rect 6825 3519 6883 3525
rect 6825 3516 6837 3519
rect 6788 3488 6837 3516
rect 6788 3476 6794 3488
rect 6825 3485 6837 3488
rect 6871 3485 6883 3519
rect 7285 3519 7343 3525
rect 7285 3516 7297 3519
rect 6825 3479 6883 3485
rect 6932 3488 7297 3516
rect 5460 3448 5488 3476
rect 4028 3420 5488 3448
rect 6564 3448 6592 3476
rect 6932 3448 6960 3488
rect 7285 3485 7297 3488
rect 7331 3485 7343 3519
rect 7285 3479 7343 3485
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3516 7987 3519
rect 8570 3516 8576 3528
rect 7975 3488 8576 3516
rect 7975 3485 7987 3488
rect 7929 3479 7987 3485
rect 6564 3420 6960 3448
rect 4028 3408 4034 3420
rect 7098 3408 7104 3460
rect 7156 3408 7162 3460
rect 7300 3448 7328 3479
rect 8570 3476 8576 3488
rect 8628 3476 8634 3528
rect 8680 3525 8708 3556
rect 9401 3553 9413 3556
rect 9447 3584 9459 3587
rect 9447 3556 10180 3584
rect 9447 3553 9459 3556
rect 9401 3547 9459 3553
rect 10152 3528 10180 3556
rect 10686 3544 10692 3596
rect 10744 3584 10750 3596
rect 10965 3587 11023 3593
rect 10965 3584 10977 3587
rect 10744 3556 10977 3584
rect 10744 3544 10750 3556
rect 10965 3553 10977 3556
rect 11011 3584 11023 3587
rect 12406 3584 12434 3692
rect 13814 3680 13820 3732
rect 13872 3720 13878 3732
rect 14737 3723 14795 3729
rect 14737 3720 14749 3723
rect 13872 3692 14749 3720
rect 13872 3680 13878 3692
rect 14737 3689 14749 3692
rect 14783 3689 14795 3723
rect 14737 3683 14795 3689
rect 12805 3655 12863 3661
rect 12805 3621 12817 3655
rect 12851 3652 12863 3655
rect 13538 3652 13544 3664
rect 12851 3624 13544 3652
rect 12851 3621 12863 3624
rect 12805 3615 12863 3621
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 14274 3612 14280 3664
rect 14332 3612 14338 3664
rect 14292 3584 14320 3612
rect 15654 3584 15660 3596
rect 11011 3556 11652 3584
rect 12406 3556 12848 3584
rect 11011 3553 11023 3556
rect 10965 3547 11023 3553
rect 8665 3519 8723 3525
rect 8665 3485 8677 3519
rect 8711 3485 8723 3519
rect 8665 3479 8723 3485
rect 9217 3519 9275 3525
rect 9217 3485 9229 3519
rect 9263 3516 9275 3519
rect 9493 3519 9551 3525
rect 9263 3488 9444 3516
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 8846 3448 8852 3460
rect 7300 3420 8852 3448
rect 8846 3408 8852 3420
rect 8904 3408 8910 3460
rect 2774 3340 2780 3392
rect 2832 3380 2838 3392
rect 3145 3383 3203 3389
rect 3145 3380 3157 3383
rect 2832 3352 3157 3380
rect 2832 3340 2838 3352
rect 3145 3349 3157 3352
rect 3191 3349 3203 3383
rect 3145 3343 3203 3349
rect 4341 3383 4399 3389
rect 4341 3349 4353 3383
rect 4387 3380 4399 3383
rect 5994 3380 6000 3392
rect 4387 3352 6000 3380
rect 4387 3349 4399 3352
rect 4341 3343 4399 3349
rect 5994 3340 6000 3352
rect 6052 3340 6058 3392
rect 6270 3340 6276 3392
rect 6328 3380 6334 3392
rect 8938 3380 8944 3392
rect 6328 3352 8944 3380
rect 6328 3340 6334 3352
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 9033 3383 9091 3389
rect 9033 3349 9045 3383
rect 9079 3380 9091 3383
rect 9306 3380 9312 3392
rect 9079 3352 9312 3380
rect 9079 3349 9091 3352
rect 9033 3343 9091 3349
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9416 3380 9444 3488
rect 9493 3485 9505 3519
rect 9539 3485 9551 3519
rect 9493 3479 9551 3485
rect 9508 3448 9536 3479
rect 9858 3476 9864 3528
rect 9916 3476 9922 3528
rect 9950 3476 9956 3528
rect 10008 3476 10014 3528
rect 10134 3476 10140 3528
rect 10192 3476 10198 3528
rect 10226 3476 10232 3528
rect 10284 3476 10290 3528
rect 10597 3519 10655 3525
rect 10597 3485 10609 3519
rect 10643 3485 10655 3519
rect 10597 3479 10655 3485
rect 9766 3448 9772 3460
rect 9508 3420 9772 3448
rect 9766 3408 9772 3420
rect 9824 3448 9830 3460
rect 10413 3451 10471 3457
rect 10413 3448 10425 3451
rect 9824 3420 10425 3448
rect 9824 3408 9830 3420
rect 10413 3417 10425 3420
rect 10459 3417 10471 3451
rect 10612 3448 10640 3479
rect 10870 3476 10876 3528
rect 10928 3476 10934 3528
rect 11146 3476 11152 3528
rect 11204 3476 11210 3528
rect 11238 3476 11244 3528
rect 11296 3476 11302 3528
rect 11514 3476 11520 3528
rect 11572 3476 11578 3528
rect 11624 3525 11652 3556
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 11790 3476 11796 3528
rect 11848 3476 11854 3528
rect 12066 3476 12072 3528
rect 12124 3476 12130 3528
rect 12820 3525 12848 3556
rect 13004 3556 14320 3584
rect 14476 3556 15660 3584
rect 13004 3525 13032 3556
rect 12345 3519 12403 3525
rect 12345 3485 12357 3519
rect 12391 3485 12403 3519
rect 12345 3479 12403 3485
rect 12805 3519 12863 3525
rect 12805 3485 12817 3519
rect 12851 3485 12863 3519
rect 12805 3479 12863 3485
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3485 13047 3519
rect 12989 3479 13047 3485
rect 11054 3448 11060 3460
rect 10612 3420 11060 3448
rect 10413 3411 10471 3417
rect 11054 3408 11060 3420
rect 11112 3448 11118 3460
rect 11808 3448 11836 3476
rect 12360 3448 12388 3479
rect 13078 3476 13084 3528
rect 13136 3476 13142 3528
rect 13173 3519 13231 3525
rect 13173 3485 13185 3519
rect 13219 3485 13231 3519
rect 13173 3479 13231 3485
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3516 13415 3519
rect 13446 3516 13452 3528
rect 13403 3488 13452 3516
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 11112 3420 12388 3448
rect 11112 3408 11118 3420
rect 10226 3380 10232 3392
rect 9416 3352 10232 3380
rect 10226 3340 10232 3352
rect 10284 3340 10290 3392
rect 10781 3383 10839 3389
rect 10781 3349 10793 3383
rect 10827 3380 10839 3383
rect 10965 3383 11023 3389
rect 10965 3380 10977 3383
rect 10827 3352 10977 3380
rect 10827 3349 10839 3352
rect 10781 3343 10839 3349
rect 10965 3349 10977 3352
rect 11011 3349 11023 3383
rect 10965 3343 11023 3349
rect 12526 3340 12532 3392
rect 12584 3340 12590 3392
rect 13096 3380 13124 3476
rect 13188 3448 13216 3479
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 14366 3525 14372 3528
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3516 13783 3519
rect 14323 3519 14372 3525
rect 14323 3518 14335 3519
rect 14322 3516 14335 3518
rect 13771 3488 14335 3516
rect 13771 3485 13783 3488
rect 13725 3479 13783 3485
rect 14323 3485 14335 3488
rect 14369 3485 14372 3519
rect 14323 3479 14372 3485
rect 14366 3476 14372 3479
rect 14424 3476 14430 3528
rect 14476 3525 14504 3556
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 14550 3476 14556 3528
rect 14608 3516 14614 3528
rect 15212 3525 15240 3556
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 14829 3519 14887 3525
rect 14829 3516 14841 3519
rect 14608 3488 14841 3516
rect 14608 3476 14614 3488
rect 14829 3485 14841 3488
rect 14875 3485 14887 3519
rect 14829 3479 14887 3485
rect 15197 3519 15255 3525
rect 15197 3485 15209 3519
rect 15243 3485 15255 3519
rect 15197 3479 15255 3485
rect 15378 3476 15384 3528
rect 15436 3516 15442 3528
rect 16114 3516 16120 3528
rect 15436 3488 16120 3516
rect 15436 3476 15442 3488
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 13630 3448 13636 3460
rect 13188 3420 13636 3448
rect 13630 3408 13636 3420
rect 13688 3408 13694 3460
rect 14093 3451 14151 3457
rect 14093 3417 14105 3451
rect 14139 3448 14151 3451
rect 14642 3448 14648 3460
rect 14139 3420 14648 3448
rect 14139 3417 14151 3420
rect 14093 3411 14151 3417
rect 14642 3408 14648 3420
rect 14700 3408 14706 3460
rect 15289 3451 15347 3457
rect 15289 3417 15301 3451
rect 15335 3448 15347 3451
rect 16574 3448 16580 3460
rect 15335 3420 16580 3448
rect 15335 3417 15347 3420
rect 15289 3411 15347 3417
rect 16574 3408 16580 3420
rect 16632 3408 16638 3460
rect 13357 3383 13415 3389
rect 13357 3380 13369 3383
rect 13096 3352 13369 3380
rect 13357 3349 13369 3352
rect 13403 3349 13415 3383
rect 13357 3343 13415 3349
rect 1104 3290 18400 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 18400 3290
rect 1104 3216 18400 3238
rect 5350 3136 5356 3188
rect 5408 3176 5414 3188
rect 5408 3148 7144 3176
rect 5408 3136 5414 3148
rect 4706 3068 4712 3120
rect 4764 3108 4770 3120
rect 6365 3111 6423 3117
rect 6365 3108 6377 3111
rect 4764 3080 6377 3108
rect 4764 3068 4770 3080
rect 6365 3077 6377 3080
rect 6411 3077 6423 3111
rect 6365 3071 6423 3077
rect 7116 3049 7144 3148
rect 7190 3136 7196 3188
rect 7248 3176 7254 3188
rect 7377 3179 7435 3185
rect 7377 3176 7389 3179
rect 7248 3148 7389 3176
rect 7248 3136 7254 3148
rect 7377 3145 7389 3148
rect 7423 3145 7435 3179
rect 7377 3139 7435 3145
rect 8938 3136 8944 3188
rect 8996 3176 9002 3188
rect 8996 3148 10088 3176
rect 8996 3136 9002 3148
rect 9677 3111 9735 3117
rect 9677 3077 9689 3111
rect 9723 3108 9735 3111
rect 9723 3080 9996 3108
rect 9723 3077 9735 3080
rect 9677 3071 9735 3077
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 7102 3043 7160 3049
rect 7102 3009 7114 3043
rect 7148 3009 7160 3043
rect 7102 3003 7160 3009
rect 5994 2932 6000 2984
rect 6052 2972 6058 2984
rect 7024 2972 7052 3003
rect 8662 3000 8668 3052
rect 8720 3040 8726 3052
rect 9033 3043 9091 3049
rect 9033 3040 9045 3043
rect 8720 3012 9045 3040
rect 8720 3000 8726 3012
rect 9033 3009 9045 3012
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3009 9275 3043
rect 9217 3003 9275 3009
rect 8570 2972 8576 2984
rect 6052 2944 6960 2972
rect 7024 2944 8576 2972
rect 6052 2932 6058 2944
rect 6086 2864 6092 2916
rect 6144 2904 6150 2916
rect 6641 2907 6699 2913
rect 6641 2904 6653 2907
rect 6144 2876 6653 2904
rect 6144 2864 6150 2876
rect 6641 2873 6653 2876
rect 6687 2873 6699 2907
rect 6641 2867 6699 2873
rect 6362 2796 6368 2848
rect 6420 2836 6426 2848
rect 6825 2839 6883 2845
rect 6825 2836 6837 2839
rect 6420 2808 6837 2836
rect 6420 2796 6426 2808
rect 6825 2805 6837 2808
rect 6871 2805 6883 2839
rect 6932 2836 6960 2944
rect 8570 2932 8576 2944
rect 8628 2932 8634 2984
rect 9232 2972 9260 3003
rect 9306 3000 9312 3052
rect 9364 3000 9370 3052
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3040 9459 3043
rect 9582 3040 9588 3052
rect 9447 3012 9588 3040
rect 9447 3009 9459 3012
rect 9401 3003 9459 3009
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 9968 3049 9996 3080
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3009 10011 3043
rect 9953 3003 10011 3009
rect 9674 2972 9680 2984
rect 9232 2944 9680 2972
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 9766 2932 9772 2984
rect 9824 2932 9830 2984
rect 10060 2972 10088 3148
rect 10134 3136 10140 3188
rect 10192 3176 10198 3188
rect 10413 3179 10471 3185
rect 10413 3176 10425 3179
rect 10192 3148 10425 3176
rect 10192 3136 10198 3148
rect 10413 3145 10425 3148
rect 10459 3145 10471 3179
rect 10413 3139 10471 3145
rect 10870 3136 10876 3188
rect 10928 3136 10934 3188
rect 12066 3136 12072 3188
rect 12124 3176 12130 3188
rect 12253 3179 12311 3185
rect 12253 3176 12265 3179
rect 12124 3148 12265 3176
rect 12124 3136 12130 3148
rect 12253 3145 12265 3148
rect 12299 3145 12311 3179
rect 12253 3139 12311 3145
rect 12526 3136 12532 3188
rect 12584 3176 12590 3188
rect 12584 3148 13400 3176
rect 12584 3136 12590 3148
rect 10594 3108 10600 3120
rect 10152 3080 10600 3108
rect 10152 3049 10180 3080
rect 10594 3068 10600 3080
rect 10652 3068 10658 3120
rect 12710 3068 12716 3120
rect 12768 3068 12774 3120
rect 12894 3068 12900 3120
rect 12952 3068 12958 3120
rect 12989 3111 13047 3117
rect 12989 3077 13001 3111
rect 13035 3108 13047 3111
rect 13265 3111 13323 3117
rect 13265 3108 13277 3111
rect 13035 3080 13277 3108
rect 13035 3077 13047 3080
rect 12989 3071 13047 3077
rect 13265 3077 13277 3080
rect 13311 3077 13323 3111
rect 13265 3071 13323 3077
rect 10137 3043 10195 3049
rect 10137 3009 10149 3043
rect 10183 3009 10195 3043
rect 10137 3003 10195 3009
rect 10226 3000 10232 3052
rect 10284 3000 10290 3052
rect 10318 3000 10324 3052
rect 10376 3000 10382 3052
rect 10410 3000 10416 3052
rect 10468 3040 10474 3052
rect 10505 3043 10563 3049
rect 10505 3040 10517 3043
rect 10468 3012 10517 3040
rect 10468 3000 10474 3012
rect 10505 3009 10517 3012
rect 10551 3009 10563 3043
rect 10505 3003 10563 3009
rect 10686 3000 10692 3052
rect 10744 3000 10750 3052
rect 10873 3043 10931 3049
rect 10873 3009 10885 3043
rect 10919 3009 10931 3043
rect 10873 3003 10931 3009
rect 10888 2972 10916 3003
rect 11606 3000 11612 3052
rect 11664 3040 11670 3052
rect 12161 3043 12219 3049
rect 12161 3040 12173 3043
rect 11664 3012 12173 3040
rect 11664 3000 11670 3012
rect 12161 3009 12173 3012
rect 12207 3009 12219 3043
rect 12345 3043 12403 3049
rect 12345 3040 12357 3043
rect 12161 3003 12219 3009
rect 12268 3012 12357 3040
rect 10060 2944 10916 2972
rect 7098 2864 7104 2916
rect 7156 2904 7162 2916
rect 7650 2904 7656 2916
rect 7156 2876 7656 2904
rect 7156 2864 7162 2876
rect 7650 2864 7656 2876
rect 7708 2904 7714 2916
rect 11882 2904 11888 2916
rect 7708 2876 11888 2904
rect 7708 2864 7714 2876
rect 11882 2864 11888 2876
rect 11940 2904 11946 2916
rect 12268 2904 12296 3012
rect 12345 3009 12357 3012
rect 12391 3009 12403 3043
rect 12345 3003 12403 3009
rect 13101 3043 13159 3049
rect 13101 3009 13113 3043
rect 13147 3040 13159 3043
rect 13372 3040 13400 3148
rect 13446 3136 13452 3188
rect 13504 3176 13510 3188
rect 15378 3176 15384 3188
rect 13504 3148 15384 3176
rect 13504 3136 13510 3148
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 13449 3043 13507 3049
rect 13449 3040 13461 3043
rect 13147 3012 13216 3040
rect 13372 3012 13461 3040
rect 13147 3009 13159 3012
rect 13101 3003 13159 3009
rect 11940 2876 12296 2904
rect 13188 2904 13216 3012
rect 13449 3009 13461 3012
rect 13495 3009 13507 3043
rect 13449 3003 13507 3009
rect 13538 3000 13544 3052
rect 13596 3000 13602 3052
rect 13262 2932 13268 2984
rect 13320 2932 13326 2984
rect 13906 2904 13912 2916
rect 13188 2876 13912 2904
rect 11940 2864 11946 2876
rect 13906 2864 13912 2876
rect 13964 2864 13970 2916
rect 11606 2836 11612 2848
rect 6932 2808 11612 2836
rect 6825 2799 6883 2805
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 12713 2839 12771 2845
rect 12713 2805 12725 2839
rect 12759 2836 12771 2839
rect 12986 2836 12992 2848
rect 12759 2808 12992 2836
rect 12759 2805 12771 2808
rect 12713 2799 12771 2805
rect 12986 2796 12992 2808
rect 13044 2796 13050 2848
rect 1104 2746 18400 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 18400 2746
rect 1104 2672 18400 2694
rect 9585 2635 9643 2641
rect 9585 2601 9597 2635
rect 9631 2632 9643 2635
rect 10226 2632 10232 2644
rect 9631 2604 10232 2632
rect 9631 2601 9643 2604
rect 9585 2595 9643 2601
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 6822 2388 6828 2440
rect 6880 2388 6886 2440
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 9490 2388 9496 2440
rect 9548 2388 9554 2440
rect 9674 2388 9680 2440
rect 9732 2388 9738 2440
rect 9766 2388 9772 2440
rect 9824 2388 9830 2440
rect 12986 2388 12992 2440
rect 13044 2428 13050 2440
rect 13633 2431 13691 2437
rect 13633 2428 13645 2431
rect 13044 2400 13645 2428
rect 13044 2388 13050 2400
rect 13633 2397 13645 2400
rect 13679 2397 13691 2431
rect 13633 2391 13691 2397
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6512 2264 6653 2292
rect 6512 2252 6518 2264
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 6641 2255 6699 2261
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 9088 2264 9321 2292
rect 9088 2252 9094 2264
rect 9309 2261 9321 2264
rect 9355 2261 9367 2295
rect 9309 2255 9367 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9953 2295 10011 2301
rect 9953 2292 9965 2295
rect 9732 2264 9965 2292
rect 9732 2252 9738 2264
rect 9953 2261 9965 2264
rect 9999 2261 10011 2295
rect 9953 2255 10011 2261
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 13817 2295 13875 2301
rect 13817 2292 13829 2295
rect 13596 2264 13829 2292
rect 13596 2252 13602 2264
rect 13817 2261 13829 2264
rect 13863 2261 13875 2295
rect 13817 2255 13875 2261
rect 1104 2202 18400 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 18400 2202
rect 1104 2128 18400 2150
<< via1 >>
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 8024 18955 8076 18964
rect 8024 18921 8033 18955
rect 8033 18921 8067 18955
rect 8067 18921 8076 18955
rect 8024 18912 8076 18921
rect 8668 18955 8720 18964
rect 8668 18921 8677 18955
rect 8677 18921 8711 18955
rect 8711 18921 8720 18955
rect 8668 18912 8720 18921
rect 9956 18955 10008 18964
rect 9956 18921 9965 18955
rect 9965 18921 9999 18955
rect 9999 18921 10008 18955
rect 9956 18912 10008 18921
rect 10600 18955 10652 18964
rect 10600 18921 10609 18955
rect 10609 18921 10643 18955
rect 10643 18921 10652 18955
rect 10600 18912 10652 18921
rect 10876 18912 10928 18964
rect 13176 18912 13228 18964
rect 7564 18708 7616 18760
rect 8484 18751 8536 18760
rect 8484 18717 8493 18751
rect 8493 18717 8527 18751
rect 8527 18717 8536 18751
rect 8484 18708 8536 18717
rect 9128 18708 9180 18760
rect 10048 18708 10100 18760
rect 11244 18708 11296 18760
rect 12348 18708 12400 18760
rect 14464 18751 14516 18760
rect 14464 18717 14473 18751
rect 14473 18717 14507 18751
rect 14507 18717 14516 18751
rect 14464 18708 14516 18717
rect 9680 18572 9732 18624
rect 13360 18615 13412 18624
rect 13360 18581 13369 18615
rect 13369 18581 13403 18615
rect 13403 18581 13412 18615
rect 13360 18572 13412 18581
rect 14740 18683 14792 18692
rect 14740 18649 14749 18683
rect 14749 18649 14783 18683
rect 14783 18649 14792 18683
rect 14740 18640 14792 18649
rect 16672 18640 16724 18692
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 7564 18411 7616 18420
rect 7564 18377 7573 18411
rect 7573 18377 7607 18411
rect 7607 18377 7616 18411
rect 7564 18368 7616 18377
rect 10048 18411 10100 18420
rect 10048 18377 10057 18411
rect 10057 18377 10091 18411
rect 10091 18377 10100 18411
rect 10048 18368 10100 18377
rect 11244 18411 11296 18420
rect 11244 18377 11253 18411
rect 11253 18377 11287 18411
rect 11287 18377 11296 18411
rect 11244 18368 11296 18377
rect 12348 18411 12400 18420
rect 12348 18377 12357 18411
rect 12357 18377 12391 18411
rect 12391 18377 12400 18411
rect 12348 18368 12400 18377
rect 7932 18275 7984 18284
rect 7932 18241 7941 18275
rect 7941 18241 7975 18275
rect 7975 18241 7984 18275
rect 7932 18232 7984 18241
rect 8116 18207 8168 18216
rect 8116 18173 8125 18207
rect 8125 18173 8159 18207
rect 8159 18173 8168 18207
rect 8116 18164 8168 18173
rect 8852 18275 8904 18284
rect 8852 18241 8861 18275
rect 8861 18241 8895 18275
rect 8895 18241 8904 18275
rect 8852 18232 8904 18241
rect 8760 18207 8812 18216
rect 8760 18173 8769 18207
rect 8769 18173 8803 18207
rect 8803 18173 8812 18207
rect 9220 18275 9272 18284
rect 9220 18241 9229 18275
rect 9229 18241 9263 18275
rect 9263 18241 9272 18275
rect 9220 18232 9272 18241
rect 8760 18164 8812 18173
rect 9128 18139 9180 18148
rect 9128 18105 9137 18139
rect 9137 18105 9171 18139
rect 9171 18105 9180 18139
rect 9128 18096 9180 18105
rect 9404 18275 9456 18284
rect 9404 18241 9413 18275
rect 9413 18241 9447 18275
rect 9447 18241 9456 18275
rect 9404 18232 9456 18241
rect 9772 18232 9824 18284
rect 10048 18232 10100 18284
rect 9680 18207 9732 18216
rect 9680 18173 9689 18207
rect 9689 18173 9723 18207
rect 9723 18173 9732 18207
rect 9680 18164 9732 18173
rect 10692 18207 10744 18216
rect 10692 18173 10701 18207
rect 10701 18173 10735 18207
rect 10735 18173 10744 18207
rect 10692 18164 10744 18173
rect 11704 18275 11756 18284
rect 11704 18241 11713 18275
rect 11713 18241 11747 18275
rect 11747 18241 11756 18275
rect 11704 18232 11756 18241
rect 16488 18300 16540 18352
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 13544 18275 13596 18284
rect 13544 18241 13553 18275
rect 13553 18241 13587 18275
rect 13587 18241 13596 18275
rect 13544 18232 13596 18241
rect 13636 18275 13688 18284
rect 13636 18241 13645 18275
rect 13645 18241 13679 18275
rect 13679 18241 13688 18275
rect 13636 18232 13688 18241
rect 16580 18232 16632 18284
rect 11796 18164 11848 18216
rect 12348 18207 12400 18216
rect 12348 18173 12357 18207
rect 12357 18173 12391 18207
rect 12391 18173 12400 18207
rect 12348 18164 12400 18173
rect 11704 18096 11756 18148
rect 13728 18096 13780 18148
rect 9680 18028 9732 18080
rect 10876 18028 10928 18080
rect 12164 18071 12216 18080
rect 12164 18037 12173 18071
rect 12173 18037 12207 18071
rect 12207 18037 12216 18071
rect 12164 18028 12216 18037
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 16764 18096 16816 18148
rect 14464 18028 14516 18080
rect 15844 18028 15896 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 8852 17824 8904 17876
rect 9404 17824 9456 17876
rect 9772 17824 9824 17876
rect 10048 17867 10100 17876
rect 10048 17833 10057 17867
rect 10057 17833 10091 17867
rect 10091 17833 10100 17867
rect 10048 17824 10100 17833
rect 10692 17867 10744 17876
rect 10692 17833 10701 17867
rect 10701 17833 10735 17867
rect 10735 17833 10744 17867
rect 10692 17824 10744 17833
rect 11520 17824 11572 17876
rect 12348 17867 12400 17876
rect 12348 17833 12357 17867
rect 12357 17833 12391 17867
rect 12391 17833 12400 17867
rect 12348 17824 12400 17833
rect 14740 17824 14792 17876
rect 16672 17867 16724 17876
rect 16672 17833 16681 17867
rect 16681 17833 16715 17867
rect 16715 17833 16724 17867
rect 16672 17824 16724 17833
rect 5724 17756 5776 17808
rect 8208 17756 8260 17808
rect 9864 17756 9916 17808
rect 12164 17756 12216 17808
rect 10600 17688 10652 17740
rect 11704 17688 11756 17740
rect 13544 17756 13596 17808
rect 14188 17756 14240 17808
rect 13360 17688 13412 17740
rect 13820 17688 13872 17740
rect 2044 17620 2096 17672
rect 8760 17620 8812 17672
rect 9220 17620 9272 17672
rect 2504 17484 2556 17536
rect 7932 17552 7984 17604
rect 9772 17552 9824 17604
rect 10876 17620 10928 17672
rect 11612 17620 11664 17672
rect 11980 17663 12032 17672
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 10416 17552 10468 17604
rect 10508 17595 10560 17604
rect 10508 17561 10517 17595
rect 10517 17561 10551 17595
rect 10551 17561 10560 17595
rect 10508 17552 10560 17561
rect 6000 17484 6052 17536
rect 8024 17484 8076 17536
rect 12992 17552 13044 17604
rect 13360 17552 13412 17604
rect 14464 17663 14516 17672
rect 14464 17629 14473 17663
rect 14473 17629 14507 17663
rect 14507 17629 14516 17663
rect 14464 17620 14516 17629
rect 15844 17620 15896 17672
rect 16580 17620 16632 17672
rect 16028 17552 16080 17604
rect 11520 17484 11572 17536
rect 14924 17484 14976 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 5724 17323 5776 17332
rect 5724 17289 5733 17323
rect 5733 17289 5767 17323
rect 5767 17289 5776 17323
rect 5724 17280 5776 17289
rect 7196 17280 7248 17332
rect 4804 17212 4856 17264
rect 3424 17076 3476 17128
rect 4068 17144 4120 17196
rect 4620 17076 4672 17128
rect 5816 17187 5868 17196
rect 5816 17153 5825 17187
rect 5825 17153 5859 17187
rect 5859 17153 5868 17187
rect 5816 17144 5868 17153
rect 6000 17144 6052 17196
rect 5540 17008 5592 17060
rect 8024 17187 8076 17196
rect 8024 17153 8033 17187
rect 8033 17153 8067 17187
rect 8067 17153 8076 17187
rect 8024 17144 8076 17153
rect 7472 17076 7524 17128
rect 8576 17187 8628 17196
rect 8576 17153 8585 17187
rect 8585 17153 8619 17187
rect 8619 17153 8628 17187
rect 8576 17144 8628 17153
rect 10416 17323 10468 17332
rect 10416 17289 10425 17323
rect 10425 17289 10459 17323
rect 10459 17289 10468 17323
rect 10416 17280 10468 17289
rect 10876 17323 10928 17332
rect 10876 17289 10885 17323
rect 10885 17289 10919 17323
rect 10919 17289 10928 17323
rect 10876 17280 10928 17289
rect 11796 17280 11848 17332
rect 12440 17280 12492 17332
rect 13636 17280 13688 17332
rect 14188 17323 14240 17332
rect 14188 17289 14197 17323
rect 14197 17289 14231 17323
rect 14231 17289 14240 17323
rect 14188 17280 14240 17289
rect 8852 17212 8904 17264
rect 8944 17187 8996 17196
rect 8944 17153 8953 17187
rect 8953 17153 8987 17187
rect 8987 17153 8996 17187
rect 10324 17212 10376 17264
rect 8944 17144 8996 17153
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 10140 17187 10192 17196
rect 10140 17153 10149 17187
rect 10149 17153 10183 17187
rect 10183 17153 10192 17187
rect 10140 17144 10192 17153
rect 9036 17008 9088 17060
rect 3792 16940 3844 16992
rect 7012 16940 7064 16992
rect 8852 16940 8904 16992
rect 9220 17119 9272 17128
rect 9220 17085 9229 17119
rect 9229 17085 9263 17119
rect 9263 17085 9272 17119
rect 9220 17076 9272 17085
rect 9772 17119 9824 17128
rect 9772 17085 9781 17119
rect 9781 17085 9815 17119
rect 9815 17085 9824 17119
rect 9772 17076 9824 17085
rect 10600 17187 10652 17196
rect 10600 17153 10609 17187
rect 10609 17153 10643 17187
rect 10643 17153 10652 17187
rect 10600 17144 10652 17153
rect 11612 17144 11664 17196
rect 11796 17187 11848 17196
rect 11796 17153 11805 17187
rect 11805 17153 11839 17187
rect 11839 17153 11848 17187
rect 11796 17144 11848 17153
rect 12256 17187 12308 17196
rect 12256 17153 12265 17187
rect 12265 17153 12299 17187
rect 12299 17153 12308 17187
rect 12256 17144 12308 17153
rect 11060 17076 11112 17128
rect 13360 17187 13412 17196
rect 13360 17153 13369 17187
rect 13369 17153 13403 17187
rect 13403 17153 13412 17187
rect 13360 17144 13412 17153
rect 16764 17255 16816 17264
rect 16764 17221 16773 17255
rect 16773 17221 16807 17255
rect 16807 17221 16816 17255
rect 16764 17212 16816 17221
rect 13728 17144 13780 17196
rect 15108 17144 15160 17196
rect 15200 17144 15252 17196
rect 11428 17008 11480 17060
rect 11796 17008 11848 17060
rect 13176 17008 13228 17060
rect 13452 17119 13504 17128
rect 13452 17085 13461 17119
rect 13461 17085 13495 17119
rect 13495 17085 13504 17119
rect 13452 17076 13504 17085
rect 13636 17076 13688 17128
rect 14096 17076 14148 17128
rect 14464 17076 14516 17128
rect 14648 17008 14700 17060
rect 16028 17008 16080 17060
rect 10416 16940 10468 16992
rect 13360 16940 13412 16992
rect 16212 16940 16264 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 8116 16736 8168 16788
rect 9864 16736 9916 16788
rect 13728 16779 13780 16788
rect 13728 16745 13737 16779
rect 13737 16745 13771 16779
rect 13771 16745 13780 16779
rect 13728 16736 13780 16745
rect 15108 16779 15160 16788
rect 15108 16745 15117 16779
rect 15117 16745 15151 16779
rect 15151 16745 15160 16779
rect 15108 16736 15160 16745
rect 3792 16600 3844 16652
rect 4068 16643 4120 16652
rect 4068 16609 4077 16643
rect 4077 16609 4111 16643
rect 4111 16609 4120 16643
rect 4068 16600 4120 16609
rect 5632 16668 5684 16720
rect 7012 16668 7064 16720
rect 2596 16532 2648 16584
rect 3424 16575 3476 16584
rect 3424 16541 3433 16575
rect 3433 16541 3467 16575
rect 3467 16541 3476 16575
rect 3424 16532 3476 16541
rect 5356 16643 5408 16652
rect 5356 16609 5365 16643
rect 5365 16609 5399 16643
rect 5399 16609 5408 16643
rect 5356 16600 5408 16609
rect 5540 16643 5592 16652
rect 5540 16609 5549 16643
rect 5549 16609 5583 16643
rect 5583 16609 5592 16643
rect 5540 16600 5592 16609
rect 8576 16668 8628 16720
rect 11796 16668 11848 16720
rect 15016 16668 15068 16720
rect 4712 16575 4764 16584
rect 4712 16541 4721 16575
rect 4721 16541 4755 16575
rect 4755 16541 4764 16575
rect 4712 16532 4764 16541
rect 4804 16575 4856 16584
rect 4804 16541 4813 16575
rect 4813 16541 4847 16575
rect 4847 16541 4856 16575
rect 4804 16532 4856 16541
rect 4988 16575 5040 16584
rect 4988 16541 4997 16575
rect 4997 16541 5031 16575
rect 5031 16541 5040 16575
rect 4988 16532 5040 16541
rect 5264 16532 5316 16584
rect 5908 16532 5960 16584
rect 6092 16575 6144 16584
rect 6092 16541 6101 16575
rect 6101 16541 6135 16575
rect 6135 16541 6144 16575
rect 6092 16532 6144 16541
rect 3056 16464 3108 16516
rect 7104 16575 7156 16584
rect 7104 16541 7113 16575
rect 7113 16541 7147 16575
rect 7147 16541 7156 16575
rect 7104 16532 7156 16541
rect 7380 16532 7432 16584
rect 7472 16575 7524 16584
rect 7472 16541 7481 16575
rect 7481 16541 7515 16575
rect 7515 16541 7524 16575
rect 7472 16532 7524 16541
rect 6460 16507 6512 16516
rect 6460 16473 6469 16507
rect 6469 16473 6503 16507
rect 6503 16473 6512 16507
rect 6460 16464 6512 16473
rect 6552 16464 6604 16516
rect 9588 16600 9640 16652
rect 8116 16575 8168 16584
rect 8116 16541 8125 16575
rect 8125 16541 8159 16575
rect 8159 16541 8168 16575
rect 8116 16532 8168 16541
rect 8760 16575 8812 16584
rect 8760 16541 8769 16575
rect 8769 16541 8803 16575
rect 8803 16541 8812 16575
rect 8760 16532 8812 16541
rect 9312 16532 9364 16584
rect 10600 16600 10652 16652
rect 9772 16532 9824 16584
rect 9956 16532 10008 16584
rect 10324 16532 10376 16584
rect 10508 16532 10560 16584
rect 12256 16600 12308 16652
rect 4988 16396 5040 16448
rect 5448 16396 5500 16448
rect 5540 16396 5592 16448
rect 6092 16396 6144 16448
rect 6828 16439 6880 16448
rect 6828 16405 6837 16439
rect 6837 16405 6871 16439
rect 6871 16405 6880 16439
rect 6828 16396 6880 16405
rect 9036 16464 9088 16516
rect 9404 16464 9456 16516
rect 11244 16532 11296 16584
rect 12900 16575 12952 16584
rect 12900 16541 12909 16575
rect 12909 16541 12943 16575
rect 12943 16541 12952 16575
rect 12900 16532 12952 16541
rect 13084 16575 13136 16584
rect 13084 16541 13093 16575
rect 13093 16541 13127 16575
rect 13127 16541 13136 16575
rect 13084 16532 13136 16541
rect 13176 16532 13228 16584
rect 13912 16600 13964 16652
rect 15844 16600 15896 16652
rect 13636 16575 13688 16584
rect 13636 16541 13645 16575
rect 13645 16541 13679 16575
rect 13679 16541 13688 16575
rect 13636 16532 13688 16541
rect 13728 16532 13780 16584
rect 12440 16464 12492 16516
rect 14832 16464 14884 16516
rect 16028 16532 16080 16584
rect 16212 16575 16264 16584
rect 16212 16541 16221 16575
rect 16221 16541 16255 16575
rect 16255 16541 16264 16575
rect 16212 16532 16264 16541
rect 16488 16575 16540 16584
rect 16488 16541 16497 16575
rect 16497 16541 16531 16575
rect 16531 16541 16540 16575
rect 16488 16532 16540 16541
rect 16580 16575 16632 16584
rect 16580 16541 16589 16575
rect 16589 16541 16623 16575
rect 16623 16541 16632 16575
rect 16580 16532 16632 16541
rect 9128 16439 9180 16448
rect 9128 16405 9137 16439
rect 9137 16405 9171 16439
rect 9171 16405 9180 16439
rect 9128 16396 9180 16405
rect 10232 16396 10284 16448
rect 13452 16439 13504 16448
rect 13452 16405 13461 16439
rect 13461 16405 13495 16439
rect 13495 16405 13504 16439
rect 13452 16396 13504 16405
rect 13728 16396 13780 16448
rect 13912 16396 13964 16448
rect 16764 16396 16816 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 2596 16056 2648 16108
rect 3056 16056 3108 16108
rect 5264 16192 5316 16244
rect 5356 16124 5408 16176
rect 5632 16235 5684 16244
rect 5632 16201 5641 16235
rect 5641 16201 5675 16235
rect 5675 16201 5684 16235
rect 5632 16192 5684 16201
rect 7840 16192 7892 16244
rect 7932 16192 7984 16244
rect 11060 16192 11112 16244
rect 14280 16192 14332 16244
rect 15844 16235 15896 16244
rect 15844 16201 15853 16235
rect 15853 16201 15887 16235
rect 15887 16201 15896 16235
rect 15844 16192 15896 16201
rect 4804 16056 4856 16108
rect 5816 16124 5868 16176
rect 6736 16167 6788 16176
rect 6736 16133 6745 16167
rect 6745 16133 6779 16167
rect 6779 16133 6788 16167
rect 6736 16124 6788 16133
rect 5080 16031 5132 16040
rect 5080 15997 5089 16031
rect 5089 15997 5123 16031
rect 5123 15997 5132 16031
rect 5080 15988 5132 15997
rect 5172 16031 5224 16040
rect 5172 15997 5181 16031
rect 5181 15997 5215 16031
rect 5215 15997 5224 16031
rect 5172 15988 5224 15997
rect 5264 16031 5316 16040
rect 5264 15997 5273 16031
rect 5273 15997 5307 16031
rect 5307 15997 5316 16031
rect 5264 15988 5316 15997
rect 6000 16056 6052 16108
rect 6828 16099 6880 16108
rect 6828 16065 6837 16099
rect 6837 16065 6871 16099
rect 6871 16065 6880 16099
rect 6828 16056 6880 16065
rect 3332 15920 3384 15972
rect 5264 15852 5316 15904
rect 5448 15920 5500 15972
rect 5724 15920 5776 15972
rect 5816 15852 5868 15904
rect 6276 15852 6328 15904
rect 6552 15895 6604 15904
rect 6552 15861 6561 15895
rect 6561 15861 6595 15895
rect 6595 15861 6604 15895
rect 6552 15852 6604 15861
rect 7104 15963 7156 15972
rect 7104 15929 7113 15963
rect 7113 15929 7147 15963
rect 7147 15929 7156 15963
rect 7104 15920 7156 15929
rect 7288 16031 7340 16040
rect 7288 15997 7297 16031
rect 7297 15997 7331 16031
rect 7331 15997 7340 16031
rect 7288 15988 7340 15997
rect 7840 16056 7892 16108
rect 8300 16056 8352 16108
rect 9036 16124 9088 16176
rect 8852 16099 8904 16108
rect 8852 16065 8861 16099
rect 8861 16065 8895 16099
rect 8895 16065 8904 16099
rect 8852 16056 8904 16065
rect 9312 16099 9364 16108
rect 9312 16065 9321 16099
rect 9321 16065 9355 16099
rect 9355 16065 9364 16099
rect 9312 16056 9364 16065
rect 9680 16056 9732 16108
rect 10140 16056 10192 16108
rect 11060 16099 11112 16108
rect 11060 16065 11069 16099
rect 11069 16065 11103 16099
rect 11103 16065 11112 16099
rect 11060 16056 11112 16065
rect 11336 16056 11388 16108
rect 12072 16167 12124 16176
rect 12072 16133 12081 16167
rect 12081 16133 12115 16167
rect 12115 16133 12124 16167
rect 12072 16124 12124 16133
rect 12256 16167 12308 16176
rect 12256 16133 12265 16167
rect 12265 16133 12299 16167
rect 12299 16133 12308 16167
rect 12256 16124 12308 16133
rect 12440 16167 12492 16176
rect 12440 16133 12449 16167
rect 12449 16133 12483 16167
rect 12483 16133 12492 16167
rect 12440 16124 12492 16133
rect 12532 16124 12584 16176
rect 13084 16167 13136 16176
rect 13084 16133 13093 16167
rect 13093 16133 13127 16167
rect 13127 16133 13136 16167
rect 13084 16124 13136 16133
rect 13636 16124 13688 16176
rect 16488 16124 16540 16176
rect 8668 15988 8720 16040
rect 9588 16031 9640 16040
rect 9588 15997 9597 16031
rect 9597 15997 9631 16031
rect 9631 15997 9640 16031
rect 9588 15988 9640 15997
rect 7564 15920 7616 15972
rect 7840 15920 7892 15972
rect 9496 15920 9548 15972
rect 8944 15852 8996 15904
rect 9128 15852 9180 15904
rect 10508 15988 10560 16040
rect 12164 16056 12216 16108
rect 13728 16056 13780 16108
rect 13820 16099 13872 16108
rect 13820 16065 13829 16099
rect 13829 16065 13863 16099
rect 13863 16065 13872 16099
rect 13820 16056 13872 16065
rect 14096 16099 14148 16108
rect 14096 16065 14105 16099
rect 14105 16065 14139 16099
rect 14139 16065 14148 16099
rect 14096 16056 14148 16065
rect 16580 16056 16632 16108
rect 17040 16056 17092 16108
rect 10784 15963 10836 15972
rect 10784 15929 10793 15963
rect 10793 15929 10827 15963
rect 10827 15929 10836 15963
rect 10784 15920 10836 15929
rect 13084 15988 13136 16040
rect 13636 16031 13688 16040
rect 13636 15997 13645 16031
rect 13645 15997 13679 16031
rect 13679 15997 13688 16031
rect 13636 15988 13688 15997
rect 13452 15920 13504 15972
rect 11060 15852 11112 15904
rect 11612 15895 11664 15904
rect 11612 15861 11621 15895
rect 11621 15861 11655 15895
rect 11655 15861 11664 15895
rect 11612 15852 11664 15861
rect 16672 15852 16724 15904
rect 17132 15852 17184 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 2964 15648 3016 15700
rect 3056 15648 3108 15700
rect 4528 15691 4580 15700
rect 4528 15657 4537 15691
rect 4537 15657 4571 15691
rect 4571 15657 4580 15691
rect 4528 15648 4580 15657
rect 6000 15648 6052 15700
rect 6552 15648 6604 15700
rect 9680 15648 9732 15700
rect 3332 15580 3384 15632
rect 3516 15512 3568 15564
rect 4620 15512 4672 15564
rect 2596 15444 2648 15496
rect 4804 15444 4856 15496
rect 6736 15580 6788 15632
rect 8024 15580 8076 15632
rect 9864 15648 9916 15700
rect 9956 15691 10008 15700
rect 9956 15657 9965 15691
rect 9965 15657 9999 15691
rect 9999 15657 10008 15691
rect 9956 15648 10008 15657
rect 11704 15648 11756 15700
rect 15752 15648 15804 15700
rect 4436 15376 4488 15428
rect 4712 15376 4764 15428
rect 6276 15512 6328 15564
rect 5540 15487 5592 15496
rect 4252 15308 4304 15360
rect 4620 15308 4672 15360
rect 5080 15376 5132 15428
rect 5172 15308 5224 15360
rect 5540 15453 5549 15487
rect 5549 15453 5583 15487
rect 5583 15453 5592 15487
rect 5540 15444 5592 15453
rect 5816 15444 5868 15496
rect 7564 15444 7616 15496
rect 7748 15487 7800 15496
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 7748 15444 7800 15453
rect 7932 15487 7984 15496
rect 7932 15453 7939 15487
rect 7939 15453 7984 15487
rect 7932 15444 7984 15453
rect 9036 15555 9088 15564
rect 9036 15521 9045 15555
rect 9045 15521 9079 15555
rect 9079 15521 9088 15555
rect 9036 15512 9088 15521
rect 8208 15487 8260 15496
rect 8208 15453 8222 15487
rect 8222 15453 8256 15487
rect 8256 15453 8260 15487
rect 8208 15444 8260 15453
rect 6092 15376 6144 15428
rect 6460 15308 6512 15360
rect 7288 15376 7340 15428
rect 8024 15419 8076 15428
rect 8024 15385 8033 15419
rect 8033 15385 8067 15419
rect 8067 15385 8076 15419
rect 8024 15376 8076 15385
rect 8760 15444 8812 15496
rect 9404 15487 9456 15496
rect 9404 15453 9413 15487
rect 9413 15453 9447 15487
rect 9447 15453 9456 15487
rect 9404 15444 9456 15453
rect 9680 15512 9732 15564
rect 17776 15580 17828 15632
rect 17224 15555 17276 15564
rect 17224 15521 17233 15555
rect 17233 15521 17267 15555
rect 17267 15521 17276 15555
rect 17224 15512 17276 15521
rect 9588 15444 9640 15496
rect 9772 15444 9824 15496
rect 12624 15444 12676 15496
rect 9312 15419 9364 15428
rect 9312 15385 9321 15419
rect 9321 15385 9355 15419
rect 9355 15385 9364 15419
rect 9312 15376 9364 15385
rect 10048 15376 10100 15428
rect 10692 15376 10744 15428
rect 12440 15376 12492 15428
rect 14924 15487 14976 15496
rect 14924 15453 14933 15487
rect 14933 15453 14967 15487
rect 14967 15453 14976 15487
rect 14924 15444 14976 15453
rect 16672 15444 16724 15496
rect 16856 15444 16908 15496
rect 17500 15487 17552 15496
rect 17500 15453 17543 15487
rect 17543 15453 17552 15487
rect 17500 15444 17552 15453
rect 8392 15351 8444 15360
rect 8392 15317 8401 15351
rect 8401 15317 8435 15351
rect 8435 15317 8444 15351
rect 8392 15308 8444 15317
rect 9864 15308 9916 15360
rect 9956 15308 10008 15360
rect 10784 15308 10836 15360
rect 12164 15308 12216 15360
rect 13176 15308 13228 15360
rect 15016 15376 15068 15428
rect 15936 15308 15988 15360
rect 16580 15308 16632 15360
rect 17592 15308 17644 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 4436 15104 4488 15156
rect 5356 15104 5408 15156
rect 7380 15104 7432 15156
rect 7932 15104 7984 15156
rect 8300 15104 8352 15156
rect 10048 15104 10100 15156
rect 2044 15011 2096 15020
rect 2044 14977 2053 15011
rect 2053 14977 2087 15011
rect 2087 14977 2096 15011
rect 2044 14968 2096 14977
rect 2412 15011 2464 15020
rect 2412 14977 2421 15011
rect 2421 14977 2455 15011
rect 2455 14977 2464 15011
rect 2412 14968 2464 14977
rect 2504 14968 2556 15020
rect 2872 14968 2924 15020
rect 3700 14968 3752 15020
rect 3976 15011 4028 15020
rect 3976 14977 3985 15011
rect 3985 14977 4019 15011
rect 4019 14977 4028 15011
rect 3976 14968 4028 14977
rect 4068 14968 4120 15020
rect 4252 15011 4304 15020
rect 4252 14977 4261 15011
rect 4261 14977 4295 15011
rect 4295 14977 4304 15011
rect 4252 14968 4304 14977
rect 2964 14943 3016 14952
rect 2964 14909 2973 14943
rect 2973 14909 3007 14943
rect 3007 14909 3016 14943
rect 2964 14900 3016 14909
rect 3240 14943 3292 14952
rect 3240 14909 3249 14943
rect 3249 14909 3283 14943
rect 3283 14909 3292 14943
rect 3240 14900 3292 14909
rect 5908 15036 5960 15088
rect 6828 15036 6880 15088
rect 8024 15036 8076 15088
rect 9404 15079 9456 15088
rect 9404 15045 9431 15079
rect 9431 15045 9456 15079
rect 9404 15036 9456 15045
rect 9588 15079 9640 15088
rect 9588 15045 9597 15079
rect 9597 15045 9631 15079
rect 9631 15045 9640 15079
rect 9588 15036 9640 15045
rect 9864 15036 9916 15088
rect 5356 14968 5408 15020
rect 7012 14968 7064 15020
rect 7380 15011 7432 15020
rect 7380 14977 7389 15011
rect 7389 14977 7423 15011
rect 7423 14977 7432 15011
rect 7380 14968 7432 14977
rect 7564 15011 7616 15020
rect 7564 14977 7573 15011
rect 7573 14977 7607 15011
rect 7607 14977 7616 15011
rect 7564 14968 7616 14977
rect 7840 14968 7892 15020
rect 7932 15011 7984 15020
rect 7932 14977 7941 15011
rect 7941 14977 7975 15011
rect 7975 14977 7984 15011
rect 7932 14968 7984 14977
rect 5540 14832 5592 14884
rect 1676 14764 1728 14816
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 2228 14764 2280 14816
rect 3240 14764 3292 14816
rect 6828 14764 6880 14816
rect 7288 14764 7340 14816
rect 7380 14764 7432 14816
rect 7564 14764 7616 14816
rect 7840 14764 7892 14816
rect 8208 14832 8260 14884
rect 10416 15011 10468 15020
rect 10416 14977 10425 15011
rect 10425 14977 10459 15011
rect 10459 14977 10468 15011
rect 10416 14968 10468 14977
rect 10692 15079 10744 15088
rect 10692 15045 10701 15079
rect 10701 15045 10735 15079
rect 10735 15045 10744 15079
rect 10692 15036 10744 15045
rect 11980 15104 12032 15156
rect 15200 15147 15252 15156
rect 15200 15113 15209 15147
rect 15209 15113 15243 15147
rect 15243 15113 15252 15147
rect 15200 15104 15252 15113
rect 15476 15104 15528 15156
rect 17040 15104 17092 15156
rect 17224 15104 17276 15156
rect 10968 15036 11020 15088
rect 12256 15036 12308 15088
rect 12808 15079 12860 15088
rect 12808 15045 12843 15079
rect 12843 15045 12860 15079
rect 12808 15036 12860 15045
rect 18052 15036 18104 15088
rect 10876 15011 10928 15020
rect 10876 14977 10885 15011
rect 10885 14977 10919 15011
rect 10919 14977 10928 15011
rect 10876 14968 10928 14977
rect 11612 14968 11664 15020
rect 12532 15011 12584 15020
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 12532 14968 12584 14977
rect 13176 14968 13228 15020
rect 13452 15011 13504 15020
rect 13452 14977 13461 15011
rect 13461 14977 13495 15011
rect 13495 14977 13504 15011
rect 13452 14968 13504 14977
rect 15752 14968 15804 15020
rect 16948 15011 17000 15020
rect 16948 14977 16957 15011
rect 16957 14977 16991 15011
rect 16991 14977 17000 15011
rect 16948 14968 17000 14977
rect 17132 14968 17184 15020
rect 17960 15011 18012 15020
rect 17960 14977 17969 15011
rect 17969 14977 18003 15011
rect 18003 14977 18012 15011
rect 17960 14968 18012 14977
rect 11428 14900 11480 14952
rect 12808 14900 12860 14952
rect 12900 14900 12952 14952
rect 12992 14943 13044 14952
rect 12992 14909 13001 14943
rect 13001 14909 13035 14943
rect 13035 14909 13044 14943
rect 12992 14900 13044 14909
rect 13084 14900 13136 14952
rect 8944 14764 8996 14816
rect 9312 14764 9364 14816
rect 13728 14900 13780 14952
rect 14556 14900 14608 14952
rect 12716 14764 12768 14816
rect 16304 14832 16356 14884
rect 17500 14832 17552 14884
rect 15476 14764 15528 14816
rect 15660 14764 15712 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 1952 14560 2004 14612
rect 2688 14560 2740 14612
rect 6460 14603 6512 14612
rect 6460 14569 6469 14603
rect 6469 14569 6503 14603
rect 6503 14569 6512 14603
rect 6460 14560 6512 14569
rect 7932 14560 7984 14612
rect 848 14492 900 14544
rect 3240 14492 3292 14544
rect 1676 14399 1728 14408
rect 1676 14365 1685 14399
rect 1685 14365 1719 14399
rect 1719 14365 1728 14399
rect 1676 14356 1728 14365
rect 2872 14424 2924 14476
rect 2412 14356 2464 14408
rect 4068 14424 4120 14476
rect 3976 14356 4028 14408
rect 4804 14424 4856 14476
rect 7564 14467 7616 14476
rect 7564 14433 7573 14467
rect 7573 14433 7607 14467
rect 7607 14433 7616 14467
rect 7564 14424 7616 14433
rect 9128 14560 9180 14612
rect 9496 14560 9548 14612
rect 9680 14560 9732 14612
rect 11520 14560 11572 14612
rect 12532 14560 12584 14612
rect 12992 14560 13044 14612
rect 8208 14492 8260 14544
rect 10968 14492 11020 14544
rect 4436 14399 4488 14408
rect 4436 14365 4445 14399
rect 4445 14365 4479 14399
rect 4479 14365 4488 14399
rect 4436 14356 4488 14365
rect 4712 14399 4764 14408
rect 4712 14365 4721 14399
rect 4721 14365 4755 14399
rect 4755 14365 4764 14399
rect 4712 14356 4764 14365
rect 4528 14263 4580 14272
rect 4528 14229 4537 14263
rect 4537 14229 4571 14263
rect 4571 14229 4580 14263
rect 4528 14220 4580 14229
rect 4712 14220 4764 14272
rect 5264 14356 5316 14408
rect 6000 14356 6052 14408
rect 5816 14288 5868 14340
rect 6552 14399 6604 14408
rect 6552 14365 6561 14399
rect 6561 14365 6595 14399
rect 6595 14365 6604 14399
rect 6552 14356 6604 14365
rect 6644 14399 6696 14408
rect 6644 14365 6653 14399
rect 6653 14365 6687 14399
rect 6687 14365 6696 14399
rect 6644 14356 6696 14365
rect 7012 14399 7064 14408
rect 7012 14365 7021 14399
rect 7021 14365 7055 14399
rect 7055 14365 7064 14399
rect 7012 14356 7064 14365
rect 6276 14288 6328 14340
rect 6828 14331 6880 14340
rect 6828 14297 6837 14331
rect 6837 14297 6871 14331
rect 6871 14297 6880 14331
rect 6828 14288 6880 14297
rect 6920 14331 6972 14340
rect 6920 14297 6929 14331
rect 6929 14297 6963 14331
rect 6963 14297 6972 14331
rect 6920 14288 6972 14297
rect 7656 14399 7708 14408
rect 7656 14365 7665 14399
rect 7665 14365 7699 14399
rect 7699 14365 7708 14399
rect 7656 14356 7708 14365
rect 8300 14356 8352 14408
rect 8024 14288 8076 14340
rect 8852 14356 8904 14408
rect 9036 14288 9088 14340
rect 6460 14220 6512 14272
rect 10508 14424 10560 14476
rect 9404 14356 9456 14408
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 9864 14356 9916 14365
rect 9956 14399 10008 14408
rect 9956 14365 9965 14399
rect 9965 14365 9999 14399
rect 9999 14365 10008 14399
rect 9956 14356 10008 14365
rect 11152 14399 11204 14408
rect 11152 14365 11161 14399
rect 11161 14365 11195 14399
rect 11195 14365 11204 14399
rect 11152 14356 11204 14365
rect 11428 14424 11480 14476
rect 11428 14331 11480 14340
rect 11428 14297 11437 14331
rect 11437 14297 11471 14331
rect 11471 14297 11480 14331
rect 11428 14288 11480 14297
rect 11520 14331 11572 14340
rect 11520 14297 11529 14331
rect 11529 14297 11563 14331
rect 11563 14297 11572 14331
rect 11520 14288 11572 14297
rect 12348 14399 12400 14408
rect 12348 14365 12357 14399
rect 12357 14365 12391 14399
rect 12391 14365 12400 14399
rect 12348 14356 12400 14365
rect 10692 14220 10744 14272
rect 12716 14467 12768 14476
rect 12716 14433 12725 14467
rect 12725 14433 12759 14467
rect 12759 14433 12768 14467
rect 12716 14424 12768 14433
rect 12900 14492 12952 14544
rect 13728 14424 13780 14476
rect 12532 14399 12584 14408
rect 12532 14365 12541 14399
rect 12541 14365 12575 14399
rect 12575 14365 12584 14399
rect 12532 14356 12584 14365
rect 12808 14356 12860 14408
rect 13912 14356 13964 14408
rect 12900 14331 12952 14340
rect 12900 14297 12909 14331
rect 12909 14297 12943 14331
rect 12943 14297 12952 14331
rect 12900 14288 12952 14297
rect 15936 14492 15988 14544
rect 16488 14492 16540 14544
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 15568 14424 15620 14476
rect 15660 14467 15712 14476
rect 15660 14433 15669 14467
rect 15669 14433 15703 14467
rect 15703 14433 15712 14467
rect 15660 14424 15712 14433
rect 15752 14467 15804 14476
rect 15752 14433 15761 14467
rect 15761 14433 15795 14467
rect 15795 14433 15804 14467
rect 15752 14424 15804 14433
rect 17684 14424 17736 14476
rect 17776 14424 17828 14476
rect 14832 14399 14884 14408
rect 14832 14365 14841 14399
rect 14841 14365 14875 14399
rect 14875 14365 14884 14399
rect 14832 14356 14884 14365
rect 15016 14356 15068 14408
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 15476 14356 15528 14408
rect 14372 14331 14424 14340
rect 14372 14297 14381 14331
rect 14381 14297 14415 14331
rect 14415 14297 14424 14331
rect 14372 14288 14424 14297
rect 14464 14331 14516 14340
rect 14464 14297 14473 14331
rect 14473 14297 14507 14331
rect 14507 14297 14516 14331
rect 14464 14288 14516 14297
rect 15476 14263 15528 14272
rect 15476 14229 15485 14263
rect 15485 14229 15519 14263
rect 15519 14229 15528 14263
rect 15476 14220 15528 14229
rect 17316 14288 17368 14340
rect 17500 14288 17552 14340
rect 17040 14220 17092 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 1584 14016 1636 14068
rect 2688 14059 2740 14068
rect 2688 14025 2697 14059
rect 2697 14025 2731 14059
rect 2731 14025 2740 14059
rect 2688 14016 2740 14025
rect 4068 14016 4120 14068
rect 4436 14016 4488 14068
rect 6736 14016 6788 14068
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 2780 13923 2832 13932
rect 2780 13889 2789 13923
rect 2789 13889 2823 13923
rect 2823 13889 2832 13923
rect 2780 13880 2832 13889
rect 3056 13923 3108 13932
rect 3056 13889 3065 13923
rect 3065 13889 3099 13923
rect 3099 13889 3108 13923
rect 3056 13880 3108 13889
rect 3240 13991 3292 14000
rect 3240 13957 3249 13991
rect 3249 13957 3283 13991
rect 3283 13957 3292 13991
rect 3240 13948 3292 13957
rect 5080 13948 5132 14000
rect 4528 13880 4580 13932
rect 5632 13948 5684 14000
rect 5724 13991 5776 14000
rect 5724 13957 5749 13991
rect 5749 13957 5776 13991
rect 5724 13948 5776 13957
rect 4068 13812 4120 13864
rect 4804 13812 4856 13864
rect 6184 13923 6236 13932
rect 6184 13889 6193 13923
rect 6193 13889 6227 13923
rect 6227 13889 6236 13923
rect 6184 13880 6236 13889
rect 6920 13923 6972 13932
rect 6920 13889 6929 13923
rect 6929 13889 6963 13923
rect 6963 13889 6972 13923
rect 6920 13880 6972 13889
rect 7104 13923 7156 13932
rect 7104 13889 7113 13923
rect 7113 13889 7147 13923
rect 7147 13889 7156 13923
rect 7104 13880 7156 13889
rect 8668 14016 8720 14068
rect 9864 14016 9916 14068
rect 11336 14016 11388 14068
rect 11428 14016 11480 14068
rect 7656 13948 7708 14000
rect 8024 13923 8076 13932
rect 8024 13889 8033 13923
rect 8033 13889 8067 13923
rect 8067 13889 8076 13923
rect 8024 13880 8076 13889
rect 8116 13880 8168 13932
rect 10600 13948 10652 14000
rect 8576 13923 8628 13932
rect 8576 13889 8585 13923
rect 8585 13889 8619 13923
rect 8619 13889 8628 13923
rect 8576 13880 8628 13889
rect 8852 13923 8904 13932
rect 8852 13889 8861 13923
rect 8861 13889 8895 13923
rect 8895 13889 8904 13923
rect 8852 13880 8904 13889
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 2320 13719 2372 13728
rect 2320 13685 2329 13719
rect 2329 13685 2363 13719
rect 2363 13685 2372 13719
rect 2320 13676 2372 13685
rect 2872 13719 2924 13728
rect 2872 13685 2881 13719
rect 2881 13685 2915 13719
rect 2915 13685 2924 13719
rect 2872 13676 2924 13685
rect 3976 13719 4028 13728
rect 3976 13685 3985 13719
rect 3985 13685 4019 13719
rect 4019 13685 4028 13719
rect 3976 13676 4028 13685
rect 5724 13719 5776 13728
rect 5724 13685 5758 13719
rect 5758 13685 5776 13719
rect 5724 13676 5776 13685
rect 6552 13812 6604 13864
rect 7840 13812 7892 13864
rect 9404 13923 9456 13932
rect 9404 13889 9413 13923
rect 9413 13889 9447 13923
rect 9447 13889 9456 13923
rect 9404 13880 9456 13889
rect 9588 13923 9640 13932
rect 9588 13889 9597 13923
rect 9597 13889 9631 13923
rect 9631 13889 9640 13923
rect 9588 13880 9640 13889
rect 9864 13880 9916 13932
rect 10784 13880 10836 13932
rect 7656 13676 7708 13728
rect 8484 13787 8536 13796
rect 8484 13753 8493 13787
rect 8493 13753 8527 13787
rect 8527 13753 8536 13787
rect 8484 13744 8536 13753
rect 8576 13744 8628 13796
rect 11704 13923 11756 13932
rect 11704 13889 11713 13923
rect 11713 13889 11747 13923
rect 11747 13889 11756 13923
rect 11704 13880 11756 13889
rect 13084 13880 13136 13932
rect 13360 13880 13412 13932
rect 13452 13880 13504 13932
rect 14372 14016 14424 14068
rect 16764 14016 16816 14068
rect 16948 14059 17000 14068
rect 16948 14025 16957 14059
rect 16957 14025 16991 14059
rect 16991 14025 17000 14059
rect 16948 14016 17000 14025
rect 17040 14059 17092 14068
rect 17040 14025 17049 14059
rect 17049 14025 17083 14059
rect 17083 14025 17092 14059
rect 17040 14016 17092 14025
rect 17500 14059 17552 14068
rect 17500 14025 17509 14059
rect 17509 14025 17543 14059
rect 17543 14025 17552 14059
rect 17500 14016 17552 14025
rect 17960 14059 18012 14068
rect 17960 14025 17969 14059
rect 17969 14025 18003 14059
rect 18003 14025 18012 14059
rect 17960 14016 18012 14025
rect 14372 13923 14424 13932
rect 14372 13889 14381 13923
rect 14381 13889 14415 13923
rect 14415 13889 14424 13923
rect 14372 13880 14424 13889
rect 12164 13855 12216 13864
rect 12164 13821 12173 13855
rect 12173 13821 12207 13855
rect 12207 13821 12216 13855
rect 12164 13812 12216 13821
rect 8760 13676 8812 13728
rect 9036 13676 9088 13728
rect 9220 13676 9272 13728
rect 9772 13719 9824 13728
rect 9772 13685 9781 13719
rect 9781 13685 9815 13719
rect 9815 13685 9824 13719
rect 9772 13676 9824 13685
rect 10692 13676 10744 13728
rect 11980 13744 12032 13796
rect 14188 13855 14240 13864
rect 14188 13821 14197 13855
rect 14197 13821 14231 13855
rect 14231 13821 14240 13855
rect 14188 13812 14240 13821
rect 14832 13948 14884 14000
rect 15476 13948 15528 14000
rect 14648 13923 14700 13932
rect 14648 13889 14657 13923
rect 14657 13889 14691 13923
rect 14691 13889 14700 13923
rect 14648 13880 14700 13889
rect 14924 13923 14976 13932
rect 14924 13889 14933 13923
rect 14933 13889 14967 13923
rect 14967 13889 14976 13923
rect 14924 13880 14976 13889
rect 15384 13880 15436 13932
rect 14832 13855 14884 13864
rect 14832 13821 14841 13855
rect 14841 13821 14875 13855
rect 14875 13821 14884 13855
rect 14832 13812 14884 13821
rect 15660 13855 15712 13864
rect 15660 13821 15669 13855
rect 15669 13821 15703 13855
rect 15703 13821 15712 13855
rect 15660 13812 15712 13821
rect 16028 13855 16080 13864
rect 16028 13821 16037 13855
rect 16037 13821 16071 13855
rect 16071 13821 16080 13855
rect 16028 13812 16080 13821
rect 16580 13880 16632 13932
rect 16764 13812 16816 13864
rect 17408 13880 17460 13932
rect 17592 13880 17644 13932
rect 17684 13880 17736 13932
rect 15108 13744 15160 13796
rect 11520 13676 11572 13728
rect 12716 13676 12768 13728
rect 14832 13676 14884 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 2872 13472 2924 13524
rect 3332 13515 3384 13524
rect 3332 13481 3341 13515
rect 3341 13481 3375 13515
rect 3375 13481 3384 13515
rect 3332 13472 3384 13481
rect 3884 13472 3936 13524
rect 4896 13472 4948 13524
rect 5448 13472 5500 13524
rect 6460 13472 6512 13524
rect 7104 13515 7156 13524
rect 7104 13481 7113 13515
rect 7113 13481 7147 13515
rect 7147 13481 7156 13515
rect 7104 13472 7156 13481
rect 7196 13472 7248 13524
rect 8024 13472 8076 13524
rect 2320 13336 2372 13388
rect 8852 13404 8904 13456
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 2504 13268 2556 13320
rect 2872 13268 2924 13320
rect 3056 13336 3108 13388
rect 3608 13336 3660 13388
rect 3148 13311 3200 13320
rect 3148 13277 3157 13311
rect 3157 13277 3191 13311
rect 3191 13277 3200 13311
rect 3148 13268 3200 13277
rect 3792 13311 3844 13320
rect 3792 13277 3801 13311
rect 3801 13277 3835 13311
rect 3835 13277 3844 13311
rect 3792 13268 3844 13277
rect 6920 13336 6972 13388
rect 10692 13472 10744 13524
rect 10876 13472 10928 13524
rect 11152 13472 11204 13524
rect 9220 13404 9272 13456
rect 10048 13404 10100 13456
rect 10968 13404 11020 13456
rect 6368 13268 6420 13320
rect 9312 13336 9364 13388
rect 12900 13404 12952 13456
rect 15292 13472 15344 13524
rect 16120 13472 16172 13524
rect 17776 13515 17828 13524
rect 17776 13481 17785 13515
rect 17785 13481 17819 13515
rect 17819 13481 17828 13515
rect 17776 13472 17828 13481
rect 1952 13132 2004 13184
rect 2872 13132 2924 13184
rect 4252 13132 4304 13184
rect 5816 13200 5868 13252
rect 7012 13200 7064 13252
rect 8576 13311 8628 13320
rect 8576 13277 8585 13311
rect 8585 13277 8619 13311
rect 8619 13277 8628 13311
rect 8576 13268 8628 13277
rect 13084 13336 13136 13388
rect 15016 13404 15068 13456
rect 17408 13404 17460 13456
rect 7932 13200 7984 13252
rect 6828 13132 6880 13184
rect 8576 13132 8628 13184
rect 8852 13200 8904 13252
rect 9312 13200 9364 13252
rect 9496 13243 9548 13252
rect 9496 13209 9505 13243
rect 9505 13209 9539 13243
rect 9539 13209 9548 13243
rect 9496 13200 9548 13209
rect 9588 13200 9640 13252
rect 10048 13311 10100 13320
rect 10048 13277 10057 13311
rect 10057 13277 10091 13311
rect 10091 13277 10100 13311
rect 10048 13268 10100 13277
rect 9680 13132 9732 13184
rect 9772 13132 9824 13184
rect 10416 13311 10468 13320
rect 10416 13277 10425 13311
rect 10425 13277 10459 13311
rect 10459 13277 10468 13311
rect 10416 13268 10468 13277
rect 10692 13268 10744 13320
rect 12992 13311 13044 13320
rect 12992 13277 13001 13311
rect 13001 13277 13035 13311
rect 13035 13277 13044 13311
rect 15752 13336 15804 13388
rect 12992 13268 13044 13277
rect 12256 13200 12308 13252
rect 12716 13132 12768 13184
rect 13820 13268 13872 13320
rect 14740 13268 14792 13320
rect 15016 13268 15068 13320
rect 14280 13200 14332 13252
rect 15660 13268 15712 13320
rect 15936 13268 15988 13320
rect 15292 13200 15344 13252
rect 13360 13132 13412 13184
rect 13728 13132 13780 13184
rect 15016 13175 15068 13184
rect 15016 13141 15025 13175
rect 15025 13141 15059 13175
rect 15059 13141 15068 13175
rect 15016 13132 15068 13141
rect 15660 13132 15712 13184
rect 16396 13132 16448 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 1676 12928 1728 12980
rect 1952 12971 2004 12980
rect 1952 12937 1961 12971
rect 1961 12937 1995 12971
rect 1995 12937 2004 12971
rect 1952 12928 2004 12937
rect 2688 12928 2740 12980
rect 3332 12928 3384 12980
rect 2872 12860 2924 12912
rect 3516 12860 3568 12912
rect 2044 12767 2096 12776
rect 2044 12733 2053 12767
rect 2053 12733 2087 12767
rect 2087 12733 2096 12767
rect 2044 12724 2096 12733
rect 2412 12724 2464 12776
rect 3056 12835 3108 12844
rect 3056 12801 3065 12835
rect 3065 12801 3099 12835
rect 3099 12801 3108 12835
rect 3056 12792 3108 12801
rect 3332 12792 3384 12844
rect 3148 12724 3200 12776
rect 3240 12724 3292 12776
rect 3884 12835 3936 12844
rect 3884 12801 3893 12835
rect 3893 12801 3927 12835
rect 3927 12801 3936 12835
rect 3884 12792 3936 12801
rect 4160 12792 4212 12844
rect 4252 12835 4304 12844
rect 4252 12801 4261 12835
rect 4261 12801 4295 12835
rect 4295 12801 4304 12835
rect 4252 12792 4304 12801
rect 5540 12928 5592 12980
rect 6368 12971 6420 12980
rect 6368 12937 6377 12971
rect 6377 12937 6411 12971
rect 6411 12937 6420 12971
rect 6368 12928 6420 12937
rect 4620 12860 4672 12912
rect 4896 12835 4948 12844
rect 4896 12801 4905 12835
rect 4905 12801 4939 12835
rect 4939 12801 4948 12835
rect 4896 12792 4948 12801
rect 5080 12835 5132 12844
rect 5080 12801 5089 12835
rect 5089 12801 5123 12835
rect 5123 12801 5132 12835
rect 5080 12792 5132 12801
rect 5908 12835 5960 12844
rect 5908 12801 5917 12835
rect 5917 12801 5951 12835
rect 5951 12801 5960 12835
rect 5908 12792 5960 12801
rect 6092 12835 6144 12844
rect 6092 12801 6101 12835
rect 6101 12801 6135 12835
rect 6135 12801 6144 12835
rect 6092 12792 6144 12801
rect 6460 12792 6512 12844
rect 6184 12767 6236 12776
rect 6184 12733 6193 12767
rect 6193 12733 6227 12767
rect 6227 12733 6236 12767
rect 6184 12724 6236 12733
rect 6736 12835 6788 12844
rect 6736 12801 6745 12835
rect 6745 12801 6779 12835
rect 6779 12801 6788 12835
rect 6736 12792 6788 12801
rect 9220 12860 9272 12912
rect 9588 12860 9640 12912
rect 9680 12860 9732 12912
rect 6920 12724 6972 12776
rect 7104 12724 7156 12776
rect 9128 12835 9180 12844
rect 9128 12801 9137 12835
rect 9137 12801 9171 12835
rect 9171 12801 9180 12835
rect 9128 12792 9180 12801
rect 9312 12792 9364 12844
rect 10416 12860 10468 12912
rect 10600 12860 10652 12912
rect 12348 12928 12400 12980
rect 12992 12928 13044 12980
rect 9680 12767 9732 12776
rect 9680 12733 9689 12767
rect 9689 12733 9723 12767
rect 9723 12733 9732 12767
rect 9680 12724 9732 12733
rect 3700 12656 3752 12708
rect 3516 12588 3568 12640
rect 3792 12588 3844 12640
rect 4620 12631 4672 12640
rect 4620 12597 4629 12631
rect 4629 12597 4663 12631
rect 4663 12597 4672 12631
rect 4620 12588 4672 12597
rect 6368 12656 6420 12708
rect 6736 12656 6788 12708
rect 10784 12835 10836 12844
rect 10784 12801 10793 12835
rect 10793 12801 10827 12835
rect 10827 12801 10836 12835
rect 10784 12792 10836 12801
rect 11612 12792 11664 12844
rect 11520 12767 11572 12776
rect 11520 12733 11529 12767
rect 11529 12733 11563 12767
rect 11563 12733 11572 12767
rect 11520 12724 11572 12733
rect 11336 12656 11388 12708
rect 11888 12835 11940 12844
rect 11888 12801 11897 12835
rect 11897 12801 11931 12835
rect 11931 12801 11940 12835
rect 11888 12792 11940 12801
rect 11980 12835 12032 12844
rect 11980 12801 11989 12835
rect 11989 12801 12023 12835
rect 12023 12801 12032 12835
rect 11980 12792 12032 12801
rect 12716 12792 12768 12844
rect 13084 12835 13136 12844
rect 13084 12801 13093 12835
rect 13093 12801 13127 12835
rect 13127 12801 13136 12835
rect 13084 12792 13136 12801
rect 13360 12792 13412 12844
rect 12256 12724 12308 12776
rect 12348 12656 12400 12708
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 14556 12860 14608 12912
rect 15016 12860 15068 12912
rect 17316 12928 17368 12980
rect 14280 12792 14332 12844
rect 14464 12792 14516 12844
rect 14740 12792 14792 12844
rect 16396 12860 16448 12912
rect 15752 12792 15804 12844
rect 16120 12835 16172 12844
rect 16120 12801 16129 12835
rect 16129 12801 16163 12835
rect 16163 12801 16172 12835
rect 16120 12792 16172 12801
rect 16304 12792 16356 12844
rect 17224 12792 17276 12844
rect 14832 12656 14884 12708
rect 15016 12699 15068 12708
rect 15016 12665 15025 12699
rect 15025 12665 15059 12699
rect 15059 12665 15068 12699
rect 15016 12656 15068 12665
rect 16396 12656 16448 12708
rect 10692 12588 10744 12640
rect 11060 12588 11112 12640
rect 11428 12588 11480 12640
rect 13176 12631 13228 12640
rect 13176 12597 13185 12631
rect 13185 12597 13219 12631
rect 13219 12597 13228 12631
rect 13176 12588 13228 12597
rect 13912 12631 13964 12640
rect 13912 12597 13921 12631
rect 13921 12597 13955 12631
rect 13955 12597 13964 12631
rect 13912 12588 13964 12597
rect 14004 12588 14056 12640
rect 14464 12588 14516 12640
rect 15844 12588 15896 12640
rect 16212 12588 16264 12640
rect 17500 12631 17552 12640
rect 17500 12597 17509 12631
rect 17509 12597 17543 12631
rect 17543 12597 17552 12631
rect 17500 12588 17552 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 2964 12384 3016 12436
rect 3884 12384 3936 12436
rect 4160 12384 4212 12436
rect 3332 12316 3384 12368
rect 4068 12316 4120 12368
rect 4620 12316 4672 12368
rect 6736 12427 6788 12436
rect 6736 12393 6745 12427
rect 6745 12393 6779 12427
rect 6779 12393 6788 12427
rect 6736 12384 6788 12393
rect 3884 12248 3936 12300
rect 4528 12248 4580 12300
rect 2964 12223 3016 12232
rect 2964 12189 2973 12223
rect 2973 12189 3007 12223
rect 3007 12189 3016 12223
rect 2964 12180 3016 12189
rect 3240 12180 3292 12232
rect 4436 12223 4488 12232
rect 4436 12189 4445 12223
rect 4445 12189 4479 12223
rect 4479 12189 4488 12223
rect 4436 12180 4488 12189
rect 5724 12359 5776 12368
rect 5724 12325 5733 12359
rect 5733 12325 5767 12359
rect 5767 12325 5776 12359
rect 5724 12316 5776 12325
rect 5908 12316 5960 12368
rect 5540 12248 5592 12300
rect 6368 12248 6420 12300
rect 7196 12316 7248 12368
rect 7748 12427 7800 12436
rect 7748 12393 7757 12427
rect 7757 12393 7791 12427
rect 7791 12393 7800 12427
rect 7748 12384 7800 12393
rect 7840 12384 7892 12436
rect 9864 12384 9916 12436
rect 10324 12384 10376 12436
rect 11520 12384 11572 12436
rect 6736 12248 6788 12300
rect 8300 12316 8352 12368
rect 8484 12316 8536 12368
rect 3424 12112 3476 12164
rect 3884 12112 3936 12164
rect 4620 12155 4672 12164
rect 4620 12121 4629 12155
rect 4629 12121 4663 12155
rect 4663 12121 4672 12155
rect 5448 12223 5500 12232
rect 5448 12189 5457 12223
rect 5457 12189 5491 12223
rect 5491 12189 5500 12223
rect 5448 12180 5500 12189
rect 7104 12180 7156 12232
rect 7196 12223 7248 12232
rect 7196 12189 7205 12223
rect 7205 12189 7239 12223
rect 7239 12189 7248 12223
rect 7196 12180 7248 12189
rect 7288 12223 7340 12232
rect 7288 12189 7297 12223
rect 7297 12189 7331 12223
rect 7331 12189 7340 12223
rect 7288 12180 7340 12189
rect 7380 12223 7432 12232
rect 7380 12189 7389 12223
rect 7389 12189 7423 12223
rect 7423 12189 7432 12223
rect 7380 12180 7432 12189
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 8760 12248 8812 12300
rect 9680 12316 9732 12368
rect 10600 12316 10652 12368
rect 7840 12180 7892 12232
rect 8024 12180 8076 12232
rect 8852 12180 8904 12232
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 9956 12248 10008 12300
rect 10232 12248 10284 12300
rect 10508 12180 10560 12232
rect 4620 12112 4672 12121
rect 2872 12044 2924 12096
rect 3516 12044 3568 12096
rect 5356 12044 5408 12096
rect 7196 12044 7248 12096
rect 7748 12044 7800 12096
rect 8576 12155 8628 12164
rect 8576 12121 8585 12155
rect 8585 12121 8619 12155
rect 8619 12121 8628 12155
rect 8576 12112 8628 12121
rect 9128 12087 9180 12096
rect 9128 12053 9137 12087
rect 9137 12053 9171 12087
rect 9171 12053 9180 12087
rect 9128 12044 9180 12053
rect 9404 12044 9456 12096
rect 10048 12112 10100 12164
rect 10876 12248 10928 12300
rect 11060 12223 11112 12232
rect 11060 12189 11069 12223
rect 11069 12189 11103 12223
rect 11103 12189 11112 12223
rect 11060 12180 11112 12189
rect 11244 12223 11296 12232
rect 11244 12189 11253 12223
rect 11253 12189 11287 12223
rect 11287 12189 11296 12223
rect 11244 12180 11296 12189
rect 11428 12291 11480 12300
rect 11428 12257 11437 12291
rect 11437 12257 11471 12291
rect 11471 12257 11480 12291
rect 11428 12248 11480 12257
rect 11704 12180 11756 12232
rect 10784 12112 10836 12164
rect 11428 12112 11480 12164
rect 13452 12384 13504 12436
rect 12348 12180 12400 12232
rect 13728 12316 13780 12368
rect 14188 12316 14240 12368
rect 14556 12316 14608 12368
rect 15200 12384 15252 12436
rect 15936 12427 15988 12436
rect 15936 12393 15945 12427
rect 15945 12393 15979 12427
rect 15979 12393 15988 12427
rect 15936 12384 15988 12393
rect 15660 12316 15712 12368
rect 13176 12223 13228 12232
rect 13176 12189 13185 12223
rect 13185 12189 13219 12223
rect 13219 12189 13228 12223
rect 13176 12180 13228 12189
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 13544 12223 13596 12232
rect 13544 12189 13553 12223
rect 13553 12189 13587 12223
rect 13587 12189 13596 12223
rect 13544 12180 13596 12189
rect 11244 12044 11296 12096
rect 11520 12044 11572 12096
rect 12348 12044 12400 12096
rect 12992 12087 13044 12096
rect 12992 12053 13001 12087
rect 13001 12053 13035 12087
rect 13035 12053 13044 12087
rect 12992 12044 13044 12053
rect 13268 12112 13320 12164
rect 16212 12248 16264 12300
rect 14372 12223 14424 12232
rect 14372 12189 14381 12223
rect 14381 12189 14415 12223
rect 14415 12189 14424 12223
rect 14372 12180 14424 12189
rect 14464 12223 14516 12232
rect 14464 12189 14473 12223
rect 14473 12189 14507 12223
rect 14507 12189 14516 12223
rect 14464 12180 14516 12189
rect 14464 12044 14516 12096
rect 14832 12180 14884 12232
rect 14648 12044 14700 12096
rect 14832 12044 14884 12096
rect 15016 12044 15068 12096
rect 17684 12223 17736 12232
rect 17684 12189 17693 12223
rect 17693 12189 17727 12223
rect 17727 12189 17736 12223
rect 17684 12180 17736 12189
rect 16396 12112 16448 12164
rect 17316 12112 17368 12164
rect 15292 12087 15344 12096
rect 15292 12053 15301 12087
rect 15301 12053 15335 12087
rect 15335 12053 15344 12087
rect 15292 12044 15344 12053
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 2964 11840 3016 11892
rect 3240 11840 3292 11892
rect 3516 11772 3568 11824
rect 4436 11840 4488 11892
rect 6460 11840 6512 11892
rect 7196 11883 7248 11892
rect 7196 11849 7205 11883
rect 7205 11849 7239 11883
rect 7239 11849 7248 11883
rect 7196 11840 7248 11849
rect 7380 11840 7432 11892
rect 5540 11772 5592 11824
rect 5908 11772 5960 11824
rect 7564 11772 7616 11824
rect 8944 11772 8996 11824
rect 10508 11840 10560 11892
rect 2596 11704 2648 11756
rect 2964 11747 3016 11756
rect 2964 11713 2973 11747
rect 2973 11713 3007 11747
rect 3007 11713 3016 11747
rect 2964 11704 3016 11713
rect 3424 11704 3476 11756
rect 3792 11747 3844 11756
rect 3792 11713 3802 11747
rect 3802 11713 3836 11747
rect 3836 11713 3844 11747
rect 3792 11704 3844 11713
rect 4068 11747 4120 11756
rect 4068 11713 4077 11747
rect 4077 11713 4111 11747
rect 4111 11713 4120 11747
rect 4068 11704 4120 11713
rect 2688 11679 2740 11688
rect 2688 11645 2697 11679
rect 2697 11645 2731 11679
rect 2731 11645 2740 11679
rect 2688 11636 2740 11645
rect 2872 11636 2924 11688
rect 4620 11704 4672 11756
rect 8024 11747 8076 11756
rect 8024 11713 8033 11747
rect 8033 11713 8067 11747
rect 8067 11713 8076 11747
rect 8024 11704 8076 11713
rect 8116 11747 8168 11756
rect 8116 11713 8125 11747
rect 8125 11713 8159 11747
rect 8159 11713 8168 11747
rect 8116 11704 8168 11713
rect 8300 11747 8352 11756
rect 8300 11713 8309 11747
rect 8309 11713 8343 11747
rect 8343 11713 8352 11747
rect 8300 11704 8352 11713
rect 8668 11704 8720 11756
rect 9312 11747 9364 11756
rect 9312 11713 9343 11747
rect 9343 11713 9364 11747
rect 9312 11704 9364 11713
rect 9404 11747 9456 11756
rect 9404 11713 9415 11747
rect 9415 11713 9449 11747
rect 9449 11713 9456 11747
rect 11796 11772 11848 11824
rect 13544 11840 13596 11892
rect 14648 11840 14700 11892
rect 9404 11704 9456 11713
rect 6000 11636 6052 11688
rect 6736 11636 6788 11688
rect 7564 11636 7616 11688
rect 9496 11636 9548 11688
rect 9680 11636 9732 11688
rect 6644 11568 6696 11620
rect 4896 11500 4948 11552
rect 6736 11500 6788 11552
rect 6920 11543 6972 11552
rect 6920 11509 6929 11543
rect 6929 11509 6963 11543
rect 6963 11509 6972 11543
rect 6920 11500 6972 11509
rect 7932 11568 7984 11620
rect 8116 11568 8168 11620
rect 8300 11568 8352 11620
rect 8484 11568 8536 11620
rect 9128 11500 9180 11552
rect 9588 11568 9640 11620
rect 9772 11568 9824 11620
rect 9680 11500 9732 11552
rect 9864 11500 9916 11552
rect 10324 11704 10376 11756
rect 12072 11704 12124 11756
rect 13728 11772 13780 11824
rect 12900 11747 12952 11756
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 12348 11636 12400 11688
rect 14096 11747 14148 11756
rect 14096 11713 14105 11747
rect 14105 11713 14139 11747
rect 14139 11713 14148 11747
rect 14096 11704 14148 11713
rect 14464 11704 14516 11756
rect 14648 11704 14700 11756
rect 13176 11636 13228 11688
rect 16764 11747 16816 11756
rect 16764 11713 16773 11747
rect 16773 11713 16807 11747
rect 16807 11713 16816 11747
rect 16764 11704 16816 11713
rect 17960 11704 18012 11756
rect 11520 11568 11572 11620
rect 12164 11568 12216 11620
rect 12532 11611 12584 11620
rect 12532 11577 12541 11611
rect 12541 11577 12575 11611
rect 12575 11577 12584 11611
rect 12532 11568 12584 11577
rect 14372 11568 14424 11620
rect 14556 11568 14608 11620
rect 15844 11568 15896 11620
rect 16948 11611 17000 11620
rect 16948 11577 16957 11611
rect 16957 11577 16991 11611
rect 16991 11577 17000 11611
rect 16948 11568 17000 11577
rect 17592 11568 17644 11620
rect 10416 11500 10468 11552
rect 10692 11500 10744 11552
rect 12256 11500 12308 11552
rect 12716 11500 12768 11552
rect 13084 11500 13136 11552
rect 13820 11500 13872 11552
rect 15016 11500 15068 11552
rect 15660 11500 15712 11552
rect 15936 11500 15988 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 3976 11296 4028 11348
rect 4712 11296 4764 11348
rect 4068 11228 4120 11280
rect 4252 11228 4304 11280
rect 2596 11135 2648 11144
rect 2596 11101 2605 11135
rect 2605 11101 2639 11135
rect 2639 11101 2648 11135
rect 2596 11092 2648 11101
rect 2688 11092 2740 11144
rect 3424 11092 3476 11144
rect 2964 11024 3016 11076
rect 3516 11067 3568 11076
rect 3516 11033 3525 11067
rect 3525 11033 3559 11067
rect 3559 11033 3568 11067
rect 4620 11092 4672 11144
rect 4804 11092 4856 11144
rect 7564 11339 7616 11348
rect 7564 11305 7573 11339
rect 7573 11305 7607 11339
rect 7607 11305 7616 11339
rect 7564 11296 7616 11305
rect 5724 11228 5776 11280
rect 6276 11271 6328 11280
rect 6276 11237 6285 11271
rect 6285 11237 6319 11271
rect 6319 11237 6328 11271
rect 6276 11228 6328 11237
rect 6736 11228 6788 11280
rect 9496 11296 9548 11348
rect 5908 11135 5960 11144
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 5908 11092 5960 11101
rect 6000 11135 6052 11144
rect 6000 11101 6009 11135
rect 6009 11101 6043 11135
rect 6043 11101 6052 11135
rect 6000 11092 6052 11101
rect 7104 11160 7156 11212
rect 7380 11160 7432 11212
rect 7748 11203 7800 11212
rect 7748 11169 7757 11203
rect 7757 11169 7791 11203
rect 7791 11169 7800 11203
rect 7748 11160 7800 11169
rect 8944 11271 8996 11280
rect 8944 11237 8953 11271
rect 8953 11237 8987 11271
rect 8987 11237 8996 11271
rect 8944 11228 8996 11237
rect 9404 11160 9456 11212
rect 10416 11339 10468 11348
rect 10416 11305 10425 11339
rect 10425 11305 10459 11339
rect 10459 11305 10468 11339
rect 10416 11296 10468 11305
rect 9956 11228 10008 11280
rect 6644 11135 6696 11144
rect 6644 11101 6653 11135
rect 6653 11101 6687 11135
rect 6687 11101 6696 11135
rect 6644 11092 6696 11101
rect 6828 11092 6880 11144
rect 6920 11135 6972 11144
rect 6920 11101 6929 11135
rect 6929 11101 6963 11135
rect 6963 11101 6972 11135
rect 6920 11092 6972 11101
rect 3516 11024 3568 11033
rect 4896 11024 4948 11076
rect 5080 11067 5132 11076
rect 5080 11033 5089 11067
rect 5089 11033 5123 11067
rect 5123 11033 5132 11067
rect 5080 11024 5132 11033
rect 5540 11067 5592 11076
rect 5540 11033 5549 11067
rect 5549 11033 5583 11067
rect 5583 11033 5592 11067
rect 5540 11024 5592 11033
rect 5816 11024 5868 11076
rect 6092 11067 6144 11076
rect 6092 11033 6101 11067
rect 6101 11033 6135 11067
rect 6135 11033 6144 11067
rect 6092 11024 6144 11033
rect 6552 11024 6604 11076
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 8024 11135 8076 11144
rect 8024 11101 8033 11135
rect 8033 11101 8067 11135
rect 8067 11101 8076 11135
rect 8024 11092 8076 11101
rect 8208 11092 8260 11144
rect 8576 11135 8628 11144
rect 8576 11101 8585 11135
rect 8585 11101 8619 11135
rect 8619 11101 8628 11135
rect 8576 11092 8628 11101
rect 8668 11092 8720 11144
rect 2136 10999 2188 11008
rect 2136 10965 2145 10999
rect 2145 10965 2179 10999
rect 2179 10965 2188 10999
rect 2136 10956 2188 10965
rect 3700 10956 3752 11008
rect 4252 10956 4304 11008
rect 6460 10956 6512 11008
rect 7748 11024 7800 11076
rect 8760 11024 8812 11076
rect 9128 11067 9180 11076
rect 9128 11033 9137 11067
rect 9137 11033 9171 11067
rect 9171 11033 9180 11067
rect 9128 11024 9180 11033
rect 9404 11024 9456 11076
rect 9588 11092 9640 11144
rect 9772 11092 9824 11144
rect 10692 11160 10744 11212
rect 11428 11296 11480 11348
rect 11796 11339 11848 11348
rect 11796 11305 11805 11339
rect 11805 11305 11839 11339
rect 11839 11305 11848 11339
rect 11796 11296 11848 11305
rect 11888 11296 11940 11348
rect 11520 11228 11572 11280
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 10876 11092 10928 11144
rect 11152 11135 11204 11144
rect 11152 11101 11162 11135
rect 11162 11101 11196 11135
rect 11196 11101 11204 11135
rect 11152 11092 11204 11101
rect 11428 11135 11480 11144
rect 11428 11101 11437 11135
rect 11437 11101 11471 11135
rect 11471 11101 11480 11135
rect 11428 11092 11480 11101
rect 12992 11296 13044 11348
rect 12348 11160 12400 11212
rect 14556 11296 14608 11348
rect 15200 11339 15252 11348
rect 15200 11305 15209 11339
rect 15209 11305 15243 11339
rect 15243 11305 15252 11339
rect 15200 11296 15252 11305
rect 17960 11339 18012 11348
rect 17960 11305 17969 11339
rect 17969 11305 18003 11339
rect 18003 11305 18012 11339
rect 17960 11296 18012 11305
rect 14464 11228 14516 11280
rect 11980 11135 12032 11144
rect 11980 11101 11989 11135
rect 11989 11101 12023 11135
rect 12023 11101 12032 11135
rect 11980 11092 12032 11101
rect 12440 11092 12492 11144
rect 12808 11092 12860 11144
rect 13820 11135 13872 11144
rect 13820 11101 13829 11135
rect 13829 11101 13863 11135
rect 13863 11101 13872 11135
rect 13820 11092 13872 11101
rect 13912 11135 13964 11144
rect 13912 11101 13921 11135
rect 13921 11101 13955 11135
rect 13955 11101 13964 11135
rect 13912 11092 13964 11101
rect 14096 11135 14148 11144
rect 14096 11101 14105 11135
rect 14105 11101 14139 11135
rect 14139 11101 14148 11135
rect 14096 11092 14148 11101
rect 14556 11160 14608 11212
rect 14740 11228 14792 11280
rect 8300 10956 8352 11008
rect 10508 10956 10560 11008
rect 10968 10956 11020 11008
rect 12624 10956 12676 11008
rect 13544 11024 13596 11076
rect 15476 11160 15528 11212
rect 15752 11160 15804 11212
rect 15016 11135 15068 11144
rect 15016 11101 15025 11135
rect 15025 11101 15059 11135
rect 15059 11101 15068 11135
rect 15016 11092 15068 11101
rect 15660 11135 15712 11144
rect 15660 11101 15669 11135
rect 15669 11101 15703 11135
rect 15703 11101 15712 11135
rect 15660 11092 15712 11101
rect 17684 11160 17736 11212
rect 15568 11024 15620 11076
rect 13636 10956 13688 11008
rect 14280 10956 14332 11008
rect 15016 10956 15068 11008
rect 15200 10956 15252 11008
rect 15476 10999 15528 11008
rect 15476 10965 15485 10999
rect 15485 10965 15519 10999
rect 15519 10965 15528 10999
rect 15476 10956 15528 10965
rect 16212 11024 16264 11076
rect 17500 11024 17552 11076
rect 16120 10956 16172 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 2872 10727 2924 10736
rect 2872 10693 2881 10727
rect 2881 10693 2915 10727
rect 2915 10693 2924 10727
rect 2872 10684 2924 10693
rect 3424 10684 3476 10736
rect 3976 10684 4028 10736
rect 4068 10684 4120 10736
rect 4712 10684 4764 10736
rect 2136 10616 2188 10668
rect 3148 10659 3200 10668
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 3240 10659 3292 10668
rect 3240 10625 3249 10659
rect 3249 10625 3283 10659
rect 3283 10625 3292 10659
rect 3240 10616 3292 10625
rect 4528 10659 4580 10668
rect 4528 10625 4537 10659
rect 4537 10625 4571 10659
rect 4571 10625 4580 10659
rect 4528 10616 4580 10625
rect 5448 10752 5500 10804
rect 5540 10752 5592 10804
rect 6920 10752 6972 10804
rect 7932 10752 7984 10804
rect 4988 10659 5040 10668
rect 4988 10625 4997 10659
rect 4997 10625 5031 10659
rect 5031 10625 5040 10659
rect 4988 10616 5040 10625
rect 5172 10659 5224 10668
rect 5172 10625 5182 10659
rect 5182 10625 5216 10659
rect 5216 10625 5224 10659
rect 5172 10616 5224 10625
rect 3792 10548 3844 10600
rect 6276 10684 6328 10736
rect 5448 10659 5500 10668
rect 5448 10625 5457 10659
rect 5457 10625 5491 10659
rect 5491 10625 5500 10659
rect 5448 10616 5500 10625
rect 6092 10616 6144 10668
rect 8300 10684 8352 10736
rect 10048 10752 10100 10804
rect 10876 10752 10928 10804
rect 7012 10616 7064 10668
rect 8208 10616 8260 10668
rect 8760 10659 8812 10668
rect 8760 10625 8769 10659
rect 8769 10625 8803 10659
rect 8803 10625 8812 10659
rect 8760 10616 8812 10625
rect 9220 10659 9272 10668
rect 9220 10625 9229 10659
rect 9229 10625 9263 10659
rect 9263 10625 9272 10659
rect 9220 10616 9272 10625
rect 9404 10659 9456 10668
rect 9404 10625 9413 10659
rect 9413 10625 9447 10659
rect 9447 10625 9456 10659
rect 9404 10616 9456 10625
rect 10600 10684 10652 10736
rect 11520 10684 11572 10736
rect 11980 10752 12032 10804
rect 12808 10752 12860 10804
rect 10048 10659 10100 10668
rect 10048 10625 10057 10659
rect 10057 10625 10091 10659
rect 10091 10625 10100 10659
rect 10048 10616 10100 10625
rect 8576 10548 8628 10600
rect 9496 10548 9548 10600
rect 9588 10548 9640 10600
rect 10232 10659 10284 10668
rect 10232 10625 10277 10659
rect 10277 10625 10284 10659
rect 10232 10616 10284 10625
rect 10876 10616 10928 10668
rect 8944 10480 8996 10532
rect 10692 10548 10744 10600
rect 11152 10659 11204 10668
rect 11152 10625 11161 10659
rect 11161 10625 11195 10659
rect 11195 10625 11204 10659
rect 11152 10616 11204 10625
rect 3056 10412 3108 10464
rect 3332 10412 3384 10464
rect 3608 10412 3660 10464
rect 3976 10412 4028 10464
rect 4804 10412 4856 10464
rect 6828 10412 6880 10464
rect 8668 10412 8720 10464
rect 8852 10455 8904 10464
rect 8852 10421 8861 10455
rect 8861 10421 8895 10455
rect 8895 10421 8904 10455
rect 10140 10480 10192 10532
rect 11980 10616 12032 10668
rect 12164 10684 12216 10736
rect 12624 10684 12676 10736
rect 13084 10684 13136 10736
rect 13820 10684 13872 10736
rect 14924 10752 14976 10804
rect 15568 10752 15620 10804
rect 17316 10752 17368 10804
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 14280 10659 14332 10668
rect 14280 10625 14289 10659
rect 14289 10625 14323 10659
rect 14323 10625 14332 10659
rect 14280 10616 14332 10625
rect 15292 10616 15344 10668
rect 15476 10659 15528 10668
rect 15476 10625 15485 10659
rect 15485 10625 15519 10659
rect 15519 10625 15528 10659
rect 15476 10616 15528 10625
rect 15568 10659 15620 10668
rect 15568 10625 15577 10659
rect 15577 10625 15611 10659
rect 15611 10625 15620 10659
rect 15568 10616 15620 10625
rect 15752 10659 15804 10668
rect 15752 10625 15761 10659
rect 15761 10625 15795 10659
rect 15795 10625 15804 10659
rect 15752 10616 15804 10625
rect 17132 10684 17184 10736
rect 17408 10684 17460 10736
rect 16028 10616 16080 10668
rect 16396 10616 16448 10668
rect 8852 10412 8904 10421
rect 9220 10412 9272 10464
rect 9772 10412 9824 10464
rect 10692 10412 10744 10464
rect 11060 10455 11112 10464
rect 11060 10421 11069 10455
rect 11069 10421 11103 10455
rect 11103 10421 11112 10455
rect 11060 10412 11112 10421
rect 12072 10548 12124 10600
rect 15200 10548 15252 10600
rect 11796 10412 11848 10464
rect 16120 10480 16172 10532
rect 17040 10591 17092 10600
rect 17040 10557 17049 10591
rect 17049 10557 17083 10591
rect 17083 10557 17092 10591
rect 17040 10548 17092 10557
rect 17592 10480 17644 10532
rect 12716 10455 12768 10464
rect 12716 10421 12725 10455
rect 12725 10421 12759 10455
rect 12759 10421 12768 10455
rect 12716 10412 12768 10421
rect 12900 10412 12952 10464
rect 13636 10412 13688 10464
rect 14096 10412 14148 10464
rect 14740 10412 14792 10464
rect 17132 10412 17184 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 2780 10208 2832 10260
rect 4252 10208 4304 10260
rect 4804 10208 4856 10260
rect 6184 10208 6236 10260
rect 6828 10251 6880 10260
rect 6828 10217 6837 10251
rect 6837 10217 6871 10251
rect 6871 10217 6880 10251
rect 6828 10208 6880 10217
rect 6920 10208 6972 10260
rect 7288 10208 7340 10260
rect 7932 10208 7984 10260
rect 3976 10140 4028 10192
rect 2412 10072 2464 10124
rect 3516 10072 3568 10124
rect 5724 10140 5776 10192
rect 6000 10140 6052 10192
rect 6276 10140 6328 10192
rect 4252 10115 4304 10124
rect 4252 10081 4261 10115
rect 4261 10081 4295 10115
rect 4295 10081 4304 10115
rect 4252 10072 4304 10081
rect 4712 10072 4764 10124
rect 2964 10047 3016 10056
rect 2964 10013 2973 10047
rect 2973 10013 3007 10047
rect 3007 10013 3016 10047
rect 2964 10004 3016 10013
rect 3056 10047 3108 10056
rect 3056 10013 3065 10047
rect 3065 10013 3099 10047
rect 3099 10013 3108 10047
rect 3056 10004 3108 10013
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 3884 9936 3936 9988
rect 4436 10004 4488 10056
rect 4804 10047 4856 10056
rect 4252 9936 4304 9988
rect 4804 10013 4808 10047
rect 4808 10013 4842 10047
rect 4842 10013 4856 10047
rect 4804 10004 4856 10013
rect 4896 10047 4948 10056
rect 4896 10013 4905 10047
rect 4905 10013 4939 10047
rect 4939 10013 4948 10047
rect 4896 10004 4948 10013
rect 5448 10072 5500 10124
rect 5816 10072 5868 10124
rect 8576 10140 8628 10192
rect 9128 10140 9180 10192
rect 9496 10208 9548 10260
rect 10600 10208 10652 10260
rect 14556 10208 14608 10260
rect 15752 10208 15804 10260
rect 16212 10251 16264 10260
rect 16212 10217 16221 10251
rect 16221 10217 16255 10251
rect 16255 10217 16264 10251
rect 16212 10208 16264 10217
rect 16304 10208 16356 10260
rect 9864 10140 9916 10192
rect 10876 10140 10928 10192
rect 10048 10072 10100 10124
rect 11520 10072 11572 10124
rect 13176 10140 13228 10192
rect 17040 10140 17092 10192
rect 5632 9936 5684 9988
rect 6828 9936 6880 9988
rect 7196 10004 7248 10056
rect 7288 10047 7340 10056
rect 7288 10013 7297 10047
rect 7297 10013 7331 10047
rect 7331 10013 7340 10047
rect 7288 10004 7340 10013
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 8760 10047 8812 10056
rect 8760 10013 8769 10047
rect 8769 10013 8803 10047
rect 8803 10013 8812 10047
rect 8760 10004 8812 10013
rect 7564 9979 7616 9988
rect 7564 9945 7573 9979
rect 7573 9945 7607 9979
rect 7607 9945 7616 9979
rect 7564 9936 7616 9945
rect 7748 9936 7800 9988
rect 9036 10004 9088 10056
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 9496 10004 9548 10056
rect 2504 9911 2556 9920
rect 2504 9877 2513 9911
rect 2513 9877 2547 9911
rect 2547 9877 2556 9911
rect 2504 9868 2556 9877
rect 3700 9868 3752 9920
rect 4712 9868 4764 9920
rect 4896 9868 4948 9920
rect 5264 9911 5316 9920
rect 5264 9877 5273 9911
rect 5273 9877 5307 9911
rect 5307 9877 5316 9911
rect 5264 9868 5316 9877
rect 5540 9868 5592 9920
rect 6000 9911 6052 9920
rect 6000 9877 6009 9911
rect 6009 9877 6043 9911
rect 6043 9877 6052 9911
rect 6000 9868 6052 9877
rect 6552 9868 6604 9920
rect 7012 9868 7064 9920
rect 7196 9868 7248 9920
rect 7288 9911 7340 9920
rect 7288 9877 7297 9911
rect 7297 9877 7331 9911
rect 7331 9877 7340 9911
rect 7288 9868 7340 9877
rect 9680 9936 9732 9988
rect 11060 10047 11112 10056
rect 11060 10013 11069 10047
rect 11069 10013 11103 10047
rect 11103 10013 11112 10047
rect 11060 10004 11112 10013
rect 11336 10004 11388 10056
rect 11704 10004 11756 10056
rect 11888 10047 11940 10056
rect 11888 10013 11897 10047
rect 11897 10013 11931 10047
rect 11931 10013 11940 10047
rect 11888 10004 11940 10013
rect 11980 10047 12032 10056
rect 11980 10013 11989 10047
rect 11989 10013 12023 10047
rect 12023 10013 12032 10047
rect 11980 10004 12032 10013
rect 11796 9936 11848 9988
rect 12072 9979 12124 9988
rect 12072 9945 12081 9979
rect 12081 9945 12115 9979
rect 12115 9945 12124 9979
rect 12072 9936 12124 9945
rect 12164 9936 12216 9988
rect 12624 10047 12676 10056
rect 12624 10013 12633 10047
rect 12633 10013 12667 10047
rect 12667 10013 12676 10047
rect 12624 10004 12676 10013
rect 12992 10072 13044 10124
rect 13084 10047 13136 10056
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 13084 10004 13136 10013
rect 14004 10072 14056 10124
rect 14556 10072 14608 10124
rect 13636 10004 13688 10056
rect 14740 10047 14792 10056
rect 14740 10013 14749 10047
rect 14749 10013 14783 10047
rect 14783 10013 14792 10047
rect 14740 10004 14792 10013
rect 15384 10047 15436 10056
rect 15384 10013 15393 10047
rect 15393 10013 15427 10047
rect 15427 10013 15436 10047
rect 15384 10004 15436 10013
rect 15476 10004 15528 10056
rect 15844 10004 15896 10056
rect 17224 10047 17276 10056
rect 17224 10013 17233 10047
rect 17233 10013 17267 10047
rect 17267 10013 17276 10047
rect 17224 10004 17276 10013
rect 14372 9979 14424 9988
rect 10232 9868 10284 9920
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 14372 9945 14381 9979
rect 14381 9945 14415 9979
rect 14415 9945 14424 9979
rect 14372 9936 14424 9945
rect 15200 9936 15252 9988
rect 16396 9979 16448 9988
rect 16396 9945 16405 9979
rect 16405 9945 16439 9979
rect 16439 9945 16448 9979
rect 16396 9936 16448 9945
rect 16948 9936 17000 9988
rect 16028 9911 16080 9920
rect 16028 9877 16037 9911
rect 16037 9877 16071 9911
rect 16071 9877 16080 9911
rect 16028 9868 16080 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 3056 9664 3108 9716
rect 3608 9664 3660 9716
rect 4620 9664 4672 9716
rect 4896 9664 4948 9716
rect 6460 9664 6512 9716
rect 6828 9664 6880 9716
rect 7932 9664 7984 9716
rect 9588 9664 9640 9716
rect 11520 9664 11572 9716
rect 11980 9664 12032 9716
rect 2228 9528 2280 9580
rect 2504 9571 2556 9580
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 2504 9528 2556 9537
rect 3700 9596 3752 9648
rect 4252 9639 4304 9648
rect 4252 9605 4261 9639
rect 4261 9605 4295 9639
rect 4295 9605 4304 9639
rect 4252 9596 4304 9605
rect 2688 9528 2740 9580
rect 2872 9571 2924 9580
rect 2872 9537 2881 9571
rect 2881 9537 2915 9571
rect 2915 9537 2924 9571
rect 2872 9528 2924 9537
rect 3056 9528 3108 9580
rect 3332 9528 3384 9580
rect 1768 9503 1820 9512
rect 1768 9469 1777 9503
rect 1777 9469 1811 9503
rect 1811 9469 1820 9503
rect 1768 9460 1820 9469
rect 2320 9460 2372 9512
rect 2412 9460 2464 9512
rect 2964 9392 3016 9444
rect 3608 9571 3660 9580
rect 3608 9537 3617 9571
rect 3617 9537 3651 9571
rect 3651 9537 3660 9571
rect 3608 9528 3660 9537
rect 5816 9639 5868 9648
rect 5816 9605 5825 9639
rect 5825 9605 5859 9639
rect 5859 9605 5868 9639
rect 5816 9596 5868 9605
rect 4620 9571 4672 9580
rect 4620 9537 4629 9571
rect 4629 9537 4663 9571
rect 4663 9537 4672 9571
rect 4620 9528 4672 9537
rect 5172 9528 5224 9580
rect 4804 9460 4856 9512
rect 4988 9503 5040 9512
rect 4988 9469 4997 9503
rect 4997 9469 5031 9503
rect 5031 9469 5040 9503
rect 4988 9460 5040 9469
rect 5080 9460 5132 9512
rect 3976 9392 4028 9444
rect 5908 9571 5960 9580
rect 5908 9537 5917 9571
rect 5917 9537 5951 9571
rect 5951 9537 5960 9571
rect 5908 9528 5960 9537
rect 6460 9528 6512 9580
rect 7012 9528 7064 9580
rect 12624 9664 12676 9716
rect 13084 9664 13136 9716
rect 13360 9664 13412 9716
rect 12440 9639 12492 9648
rect 12440 9605 12449 9639
rect 12449 9605 12483 9639
rect 12483 9605 12492 9639
rect 12440 9596 12492 9605
rect 12532 9639 12584 9648
rect 12532 9605 12541 9639
rect 12541 9605 12575 9639
rect 12575 9605 12584 9639
rect 12532 9596 12584 9605
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 7288 9571 7340 9580
rect 7288 9537 7297 9571
rect 7297 9537 7331 9571
rect 7331 9537 7340 9571
rect 7288 9528 7340 9537
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 7932 9528 7984 9580
rect 9680 9528 9732 9580
rect 10048 9528 10100 9580
rect 10968 9528 11020 9580
rect 12072 9528 12124 9580
rect 12256 9571 12308 9580
rect 12256 9537 12265 9571
rect 12265 9537 12299 9571
rect 12299 9537 12308 9571
rect 12256 9528 12308 9537
rect 1676 9324 1728 9376
rect 3332 9324 3384 9376
rect 3516 9324 3568 9376
rect 4988 9324 5040 9376
rect 5540 9324 5592 9376
rect 6460 9324 6512 9376
rect 7012 9435 7064 9444
rect 7012 9401 7021 9435
rect 7021 9401 7055 9435
rect 7055 9401 7064 9435
rect 7012 9392 7064 9401
rect 7656 9503 7708 9512
rect 7656 9469 7665 9503
rect 7665 9469 7699 9503
rect 7699 9469 7708 9503
rect 7656 9460 7708 9469
rect 10784 9460 10836 9512
rect 11704 9460 11756 9512
rect 12532 9460 12584 9512
rect 13360 9528 13412 9580
rect 14004 9571 14056 9586
rect 14004 9537 14005 9571
rect 14005 9537 14039 9571
rect 14039 9537 14056 9571
rect 14004 9534 14056 9537
rect 14464 9664 14516 9716
rect 14556 9664 14608 9716
rect 16120 9639 16172 9648
rect 16120 9605 16129 9639
rect 16129 9605 16163 9639
rect 16163 9605 16172 9639
rect 16120 9596 16172 9605
rect 12716 9460 12768 9512
rect 14280 9571 14332 9580
rect 14280 9537 14289 9571
rect 14289 9537 14323 9571
rect 14323 9537 14332 9571
rect 14280 9528 14332 9537
rect 14372 9571 14424 9580
rect 14372 9537 14381 9571
rect 14381 9537 14415 9571
rect 14415 9537 14424 9571
rect 14372 9528 14424 9537
rect 14556 9528 14608 9580
rect 14648 9571 14700 9580
rect 14648 9537 14657 9571
rect 14657 9537 14691 9571
rect 14691 9537 14700 9571
rect 14648 9528 14700 9537
rect 14740 9571 14792 9580
rect 14740 9537 14749 9571
rect 14749 9537 14783 9571
rect 14783 9537 14792 9571
rect 14740 9528 14792 9537
rect 14924 9528 14976 9580
rect 9036 9392 9088 9444
rect 9864 9392 9916 9444
rect 6828 9324 6880 9376
rect 7380 9324 7432 9376
rect 8116 9324 8168 9376
rect 10048 9324 10100 9376
rect 11060 9324 11112 9376
rect 11612 9324 11664 9376
rect 11796 9324 11848 9376
rect 12072 9324 12124 9376
rect 13084 9392 13136 9444
rect 12716 9324 12768 9376
rect 12900 9324 12952 9376
rect 13728 9367 13780 9376
rect 13728 9333 13737 9367
rect 13737 9333 13771 9367
rect 13771 9333 13780 9367
rect 13728 9324 13780 9333
rect 15016 9460 15068 9512
rect 16672 9571 16724 9580
rect 16672 9537 16681 9571
rect 16681 9537 16715 9571
rect 16715 9537 16724 9571
rect 16672 9528 16724 9537
rect 17684 9571 17736 9580
rect 17684 9537 17693 9571
rect 17693 9537 17727 9571
rect 17727 9537 17736 9571
rect 17684 9528 17736 9537
rect 15844 9460 15896 9512
rect 15936 9460 15988 9512
rect 14464 9392 14516 9444
rect 15200 9392 15252 9444
rect 15384 9324 15436 9376
rect 16396 9367 16448 9376
rect 16396 9333 16405 9367
rect 16405 9333 16439 9367
rect 16439 9333 16448 9367
rect 16396 9324 16448 9333
rect 17040 9324 17092 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 2688 9120 2740 9172
rect 2964 9120 3016 9172
rect 2412 9052 2464 9104
rect 1676 8959 1728 8968
rect 1676 8925 1685 8959
rect 1685 8925 1719 8959
rect 1719 8925 1728 8959
rect 1676 8916 1728 8925
rect 1768 8916 1820 8968
rect 2504 8959 2556 8968
rect 2504 8925 2513 8959
rect 2513 8925 2547 8959
rect 2547 8925 2556 8959
rect 2504 8916 2556 8925
rect 2872 8916 2924 8968
rect 4436 9120 4488 9172
rect 7656 9120 7708 9172
rect 9496 9163 9548 9172
rect 9496 9129 9505 9163
rect 9505 9129 9539 9163
rect 9539 9129 9548 9163
rect 9496 9120 9548 9129
rect 11612 9120 11664 9172
rect 14464 9120 14516 9172
rect 16856 9120 16908 9172
rect 3792 9095 3844 9104
rect 3792 9061 3801 9095
rect 3801 9061 3835 9095
rect 3835 9061 3844 9095
rect 3792 9052 3844 9061
rect 3884 9052 3936 9104
rect 5080 9052 5132 9104
rect 6000 9052 6052 9104
rect 7104 9052 7156 9104
rect 8024 9052 8076 9104
rect 9036 9052 9088 9104
rect 11796 9052 11848 9104
rect 12716 9052 12768 9104
rect 13636 9052 13688 9104
rect 14004 9052 14056 9104
rect 15292 9052 15344 9104
rect 15936 9052 15988 9104
rect 3792 8916 3844 8968
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 4252 8959 4304 8968
rect 4252 8925 4261 8959
rect 4261 8925 4295 8959
rect 4295 8925 4304 8959
rect 4252 8916 4304 8925
rect 4896 8916 4948 8968
rect 2780 8891 2832 8900
rect 2780 8857 2789 8891
rect 2789 8857 2823 8891
rect 2823 8857 2832 8891
rect 2780 8848 2832 8857
rect 3056 8891 3108 8900
rect 3056 8857 3065 8891
rect 3065 8857 3099 8891
rect 3099 8857 3108 8891
rect 3056 8848 3108 8857
rect 5540 8848 5592 8900
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 7472 8984 7524 9036
rect 6920 8916 6972 8968
rect 8116 8959 8168 8968
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 8116 8916 8168 8925
rect 9680 8984 9732 9036
rect 9312 8916 9364 8968
rect 10876 8984 10928 9036
rect 9864 8959 9916 8968
rect 9864 8925 9873 8959
rect 9873 8925 9907 8959
rect 9907 8925 9916 8959
rect 9864 8916 9916 8925
rect 9956 8916 10008 8968
rect 7012 8848 7064 8900
rect 1032 8780 1084 8832
rect 3148 8780 3200 8832
rect 4620 8780 4672 8832
rect 4804 8780 4856 8832
rect 6828 8780 6880 8832
rect 7932 8891 7984 8900
rect 7932 8857 7941 8891
rect 7941 8857 7975 8891
rect 7975 8857 7984 8891
rect 7932 8848 7984 8857
rect 10416 8916 10468 8968
rect 10692 8916 10744 8968
rect 11336 8916 11388 8968
rect 14280 8984 14332 9036
rect 11704 8848 11756 8900
rect 12256 8959 12308 8968
rect 12256 8925 12265 8959
rect 12265 8925 12299 8959
rect 12299 8925 12308 8959
rect 12256 8916 12308 8925
rect 14464 8959 14516 8968
rect 14464 8925 14473 8959
rect 14473 8925 14507 8959
rect 14507 8925 14516 8959
rect 14464 8916 14516 8925
rect 14740 8959 14792 8968
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 14740 8916 14792 8925
rect 14924 8916 14976 8968
rect 8668 8780 8720 8832
rect 9588 8780 9640 8832
rect 11152 8780 11204 8832
rect 12532 8780 12584 8832
rect 13084 8780 13136 8832
rect 14188 8823 14240 8832
rect 14188 8789 14197 8823
rect 14197 8789 14231 8823
rect 14231 8789 14240 8823
rect 14188 8780 14240 8789
rect 14372 8780 14424 8832
rect 15660 8916 15712 8968
rect 16120 8959 16172 8968
rect 16120 8925 16129 8959
rect 16129 8925 16163 8959
rect 16163 8925 16172 8959
rect 16120 8916 16172 8925
rect 16212 8916 16264 8968
rect 16396 8916 16448 8968
rect 17040 8959 17092 8968
rect 17040 8925 17049 8959
rect 17049 8925 17083 8959
rect 17083 8925 17092 8959
rect 17040 8916 17092 8925
rect 17408 8959 17460 8968
rect 17408 8925 17417 8959
rect 17417 8925 17451 8959
rect 17451 8925 17460 8959
rect 17408 8916 17460 8925
rect 15660 8823 15712 8832
rect 15660 8789 15669 8823
rect 15669 8789 15703 8823
rect 15703 8789 15712 8823
rect 15660 8780 15712 8789
rect 15936 8823 15988 8832
rect 15936 8789 15945 8823
rect 15945 8789 15979 8823
rect 15979 8789 15988 8823
rect 15936 8780 15988 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 4068 8619 4120 8628
rect 4068 8585 4077 8619
rect 4077 8585 4111 8619
rect 4111 8585 4120 8619
rect 4068 8576 4120 8585
rect 4252 8576 4304 8628
rect 5724 8508 5776 8560
rect 5816 8551 5868 8560
rect 5816 8517 5825 8551
rect 5825 8517 5859 8551
rect 5859 8517 5868 8551
rect 5816 8508 5868 8517
rect 6000 8551 6052 8560
rect 6000 8517 6009 8551
rect 6009 8517 6043 8551
rect 6043 8517 6052 8551
rect 6000 8508 6052 8517
rect 4620 8440 4672 8492
rect 5172 8440 5224 8492
rect 5908 8372 5960 8424
rect 6092 8372 6144 8424
rect 6184 8347 6236 8356
rect 6184 8313 6193 8347
rect 6193 8313 6227 8347
rect 6227 8313 6236 8347
rect 6184 8304 6236 8313
rect 3976 8236 4028 8288
rect 4804 8236 4856 8288
rect 6920 8508 6972 8560
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 7012 8440 7064 8492
rect 6644 8415 6696 8424
rect 6644 8381 6653 8415
rect 6653 8381 6687 8415
rect 6687 8381 6696 8415
rect 6644 8372 6696 8381
rect 7104 8415 7156 8424
rect 7104 8381 7113 8415
rect 7113 8381 7147 8415
rect 7147 8381 7156 8415
rect 7104 8372 7156 8381
rect 7288 8415 7340 8424
rect 7288 8381 7297 8415
rect 7297 8381 7331 8415
rect 7331 8381 7340 8415
rect 7288 8372 7340 8381
rect 8484 8508 8536 8560
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 7748 8440 7800 8492
rect 7932 8440 7984 8492
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 8576 8483 8628 8492
rect 8576 8449 8585 8483
rect 8585 8449 8619 8483
rect 8619 8449 8628 8483
rect 8576 8440 8628 8449
rect 8668 8483 8720 8492
rect 8668 8449 8677 8483
rect 8677 8449 8711 8483
rect 8711 8449 8720 8483
rect 8668 8440 8720 8449
rect 8852 8483 8904 8492
rect 8852 8449 8861 8483
rect 8861 8449 8895 8483
rect 8895 8449 8904 8483
rect 8852 8440 8904 8449
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 9220 8483 9272 8492
rect 9220 8449 9229 8483
rect 9229 8449 9263 8483
rect 9263 8449 9272 8483
rect 9220 8440 9272 8449
rect 9956 8508 10008 8560
rect 11336 8576 11388 8628
rect 13268 8576 13320 8628
rect 13636 8576 13688 8628
rect 14464 8619 14516 8628
rect 14464 8585 14473 8619
rect 14473 8585 14507 8619
rect 14507 8585 14516 8619
rect 14464 8576 14516 8585
rect 14740 8576 14792 8628
rect 9496 8440 9548 8492
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 10416 8483 10468 8492
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 10692 8440 10744 8492
rect 11060 8483 11112 8492
rect 11060 8449 11069 8483
rect 11069 8449 11103 8483
rect 11103 8449 11112 8483
rect 11060 8440 11112 8449
rect 11152 8483 11204 8492
rect 11152 8449 11161 8483
rect 11161 8449 11195 8483
rect 11195 8449 11204 8483
rect 11152 8440 11204 8449
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 12256 8508 12308 8560
rect 12808 8551 12860 8560
rect 12808 8517 12817 8551
rect 12817 8517 12851 8551
rect 12851 8517 12860 8551
rect 12808 8508 12860 8517
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 12440 8440 12492 8492
rect 13636 8440 13688 8492
rect 13728 8483 13780 8492
rect 13728 8449 13737 8483
rect 13737 8449 13771 8483
rect 13771 8449 13780 8483
rect 14372 8508 14424 8560
rect 15476 8576 15528 8628
rect 16120 8576 16172 8628
rect 13728 8440 13780 8449
rect 7472 8304 7524 8356
rect 8024 8304 8076 8356
rect 8116 8236 8168 8288
rect 9588 8304 9640 8356
rect 9680 8347 9732 8356
rect 9680 8313 9689 8347
rect 9689 8313 9723 8347
rect 9723 8313 9732 8347
rect 9680 8304 9732 8313
rect 9772 8347 9824 8356
rect 9772 8313 9781 8347
rect 9781 8313 9815 8347
rect 9815 8313 9824 8347
rect 9772 8304 9824 8313
rect 10508 8304 10560 8356
rect 13268 8372 13320 8424
rect 14004 8415 14056 8424
rect 14004 8381 14013 8415
rect 14013 8381 14047 8415
rect 14047 8381 14056 8415
rect 14004 8372 14056 8381
rect 14372 8372 14424 8424
rect 14832 8483 14884 8492
rect 14832 8449 14841 8483
rect 14841 8449 14875 8483
rect 14875 8449 14884 8483
rect 14832 8440 14884 8449
rect 15936 8508 15988 8560
rect 15200 8483 15252 8492
rect 15200 8449 15209 8483
rect 15209 8449 15243 8483
rect 15243 8449 15252 8483
rect 15200 8440 15252 8449
rect 15292 8483 15344 8492
rect 15292 8449 15301 8483
rect 15301 8449 15335 8483
rect 15335 8449 15344 8483
rect 15292 8440 15344 8449
rect 15752 8440 15804 8492
rect 15844 8483 15896 8492
rect 15844 8449 15853 8483
rect 15853 8449 15887 8483
rect 15887 8449 15896 8483
rect 15844 8440 15896 8449
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 16580 8508 16632 8560
rect 16488 8483 16540 8492
rect 16488 8449 16497 8483
rect 16497 8449 16531 8483
rect 16531 8449 16540 8483
rect 16488 8440 16540 8449
rect 17040 8508 17092 8560
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 13360 8304 13412 8356
rect 14648 8304 14700 8356
rect 9496 8236 9548 8288
rect 10692 8236 10744 8288
rect 12164 8236 12216 8288
rect 12624 8236 12676 8288
rect 13728 8236 13780 8288
rect 13912 8236 13964 8288
rect 14740 8236 14792 8288
rect 15752 8236 15804 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 3608 8032 3660 8084
rect 6552 8032 6604 8084
rect 6828 8032 6880 8084
rect 4344 7964 4396 8016
rect 3516 7896 3568 7948
rect 5632 7964 5684 8016
rect 6092 7964 6144 8016
rect 6644 7896 6696 7948
rect 7380 8032 7432 8084
rect 8208 8032 8260 8084
rect 10508 8032 10560 8084
rect 10600 8032 10652 8084
rect 7564 7964 7616 8016
rect 9496 7964 9548 8016
rect 9588 7964 9640 8016
rect 11520 7964 11572 8016
rect 3332 7828 3384 7880
rect 3424 7828 3476 7880
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 4528 7828 4580 7880
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 3056 7803 3108 7812
rect 3056 7769 3065 7803
rect 3065 7769 3099 7803
rect 3099 7769 3108 7803
rect 4804 7828 4856 7880
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 3056 7760 3108 7769
rect 4528 7692 4580 7744
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 6000 7871 6052 7880
rect 6000 7837 6007 7871
rect 6007 7837 6052 7871
rect 6000 7828 6052 7837
rect 6276 7871 6328 7880
rect 6276 7837 6290 7871
rect 6290 7837 6324 7871
rect 6324 7837 6328 7871
rect 6276 7828 6328 7837
rect 5908 7692 5960 7744
rect 6000 7692 6052 7744
rect 7288 7871 7340 7880
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 9680 7896 9732 7948
rect 7840 7828 7892 7880
rect 8300 7828 8352 7880
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 9312 7828 9364 7837
rect 10508 7896 10560 7948
rect 9864 7871 9916 7880
rect 9864 7837 9868 7871
rect 9868 7837 9902 7871
rect 9902 7837 9916 7871
rect 9864 7828 9916 7837
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 6368 7692 6420 7744
rect 6920 7692 6972 7744
rect 7288 7692 7340 7744
rect 9496 7692 9548 7744
rect 9680 7735 9732 7744
rect 9680 7701 9689 7735
rect 9689 7701 9723 7735
rect 9723 7701 9732 7735
rect 9680 7692 9732 7701
rect 9956 7803 10008 7812
rect 9956 7769 9965 7803
rect 9965 7769 9999 7803
rect 9999 7769 10008 7803
rect 9956 7760 10008 7769
rect 10232 7828 10284 7880
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 11244 7871 11296 7880
rect 11244 7837 11253 7871
rect 11253 7837 11287 7871
rect 11287 7837 11296 7871
rect 11244 7828 11296 7837
rect 11336 7871 11388 7880
rect 11336 7837 11345 7871
rect 11345 7837 11379 7871
rect 11379 7837 11388 7871
rect 11336 7828 11388 7837
rect 11520 7871 11572 7880
rect 11520 7837 11529 7871
rect 11529 7837 11563 7871
rect 11563 7837 11572 7871
rect 11520 7828 11572 7837
rect 12072 7964 12124 8016
rect 12440 7964 12492 8016
rect 13176 7964 13228 8016
rect 13728 8032 13780 8084
rect 14188 8075 14240 8084
rect 14188 8041 14197 8075
rect 14197 8041 14231 8075
rect 14231 8041 14240 8075
rect 14188 8032 14240 8041
rect 15660 8032 15712 8084
rect 16120 8032 16172 8084
rect 15292 7964 15344 8016
rect 15752 7964 15804 8016
rect 12164 7896 12216 7948
rect 11980 7871 12032 7880
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12256 7828 12308 7837
rect 12624 7828 12676 7880
rect 13636 7896 13688 7948
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 14096 7871 14148 7880
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 15476 7828 15528 7880
rect 16212 7828 16264 7880
rect 10968 7692 11020 7744
rect 14648 7760 14700 7812
rect 12716 7692 12768 7744
rect 13176 7692 13228 7744
rect 15292 7692 15344 7744
rect 15844 7692 15896 7744
rect 17960 7735 18012 7744
rect 17960 7701 17969 7735
rect 17969 7701 18003 7735
rect 18003 7701 18012 7735
rect 17960 7692 18012 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 3240 7488 3292 7540
rect 3424 7352 3476 7404
rect 3516 7395 3568 7404
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 3884 7352 3936 7404
rect 4068 7352 4120 7404
rect 5356 7420 5408 7472
rect 3240 7284 3292 7336
rect 4712 7352 4764 7404
rect 6276 7488 6328 7540
rect 6552 7488 6604 7540
rect 6920 7488 6972 7540
rect 7380 7488 7432 7540
rect 7840 7488 7892 7540
rect 9680 7488 9732 7540
rect 9864 7488 9916 7540
rect 11244 7488 11296 7540
rect 12256 7488 12308 7540
rect 6000 7420 6052 7472
rect 7288 7420 7340 7472
rect 5356 7327 5408 7336
rect 5356 7293 5365 7327
rect 5365 7293 5399 7327
rect 5399 7293 5408 7327
rect 5356 7284 5408 7293
rect 3148 7216 3200 7268
rect 3516 7216 3568 7268
rect 5540 7327 5592 7336
rect 5540 7293 5549 7327
rect 5549 7293 5583 7327
rect 5583 7293 5592 7327
rect 5540 7284 5592 7293
rect 6552 7352 6604 7404
rect 7012 7352 7064 7404
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 7748 7395 7800 7404
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 9588 7420 9640 7472
rect 9496 7395 9548 7404
rect 9496 7361 9505 7395
rect 9505 7361 9539 7395
rect 9539 7361 9548 7395
rect 9496 7352 9548 7361
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 10324 7395 10376 7404
rect 10324 7361 10333 7395
rect 10333 7361 10367 7395
rect 10367 7361 10376 7395
rect 10324 7352 10376 7361
rect 7840 7284 7892 7336
rect 9036 7327 9088 7336
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 7012 7216 7064 7268
rect 10048 7284 10100 7336
rect 10692 7327 10744 7336
rect 10692 7293 10701 7327
rect 10701 7293 10735 7327
rect 10735 7293 10744 7327
rect 10692 7284 10744 7293
rect 10968 7395 11020 7404
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 11520 7420 11572 7472
rect 14096 7488 14148 7540
rect 15108 7531 15160 7540
rect 15108 7497 15117 7531
rect 15117 7497 15151 7531
rect 15151 7497 15160 7531
rect 15108 7488 15160 7497
rect 11244 7352 11296 7404
rect 11796 7395 11848 7404
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 11796 7352 11848 7361
rect 11980 7352 12032 7404
rect 12256 7352 12308 7404
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 12440 7352 12492 7361
rect 12624 7395 12676 7404
rect 12624 7361 12633 7395
rect 12633 7361 12667 7395
rect 12667 7361 12676 7395
rect 12624 7352 12676 7361
rect 14648 7420 14700 7472
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 12992 7352 13044 7361
rect 13176 7352 13228 7404
rect 13544 7395 13596 7404
rect 13544 7361 13553 7395
rect 13553 7361 13587 7395
rect 13587 7361 13596 7395
rect 13544 7352 13596 7361
rect 13636 7352 13688 7404
rect 11152 7284 11204 7336
rect 12808 7327 12860 7336
rect 12808 7293 12817 7327
rect 12817 7293 12851 7327
rect 12851 7293 12860 7327
rect 12808 7284 12860 7293
rect 13912 7395 13964 7404
rect 13912 7361 13921 7395
rect 13921 7361 13955 7395
rect 13955 7361 13964 7395
rect 13912 7352 13964 7361
rect 14004 7352 14056 7404
rect 14188 7352 14240 7404
rect 15292 7395 15344 7404
rect 15292 7361 15301 7395
rect 15301 7361 15335 7395
rect 15335 7361 15344 7395
rect 15292 7352 15344 7361
rect 15752 7395 15804 7404
rect 15752 7361 15761 7395
rect 15761 7361 15795 7395
rect 15795 7361 15804 7395
rect 15752 7352 15804 7361
rect 16212 7395 16264 7404
rect 16212 7361 16221 7395
rect 16221 7361 16255 7395
rect 16255 7361 16264 7395
rect 16212 7352 16264 7361
rect 16948 7352 17000 7404
rect 2872 7191 2924 7200
rect 2872 7157 2881 7191
rect 2881 7157 2915 7191
rect 2915 7157 2924 7191
rect 2872 7148 2924 7157
rect 3700 7148 3752 7200
rect 3792 7148 3844 7200
rect 4344 7191 4396 7200
rect 4344 7157 4353 7191
rect 4353 7157 4387 7191
rect 4387 7157 4396 7191
rect 4344 7148 4396 7157
rect 5632 7148 5684 7200
rect 6460 7148 6512 7200
rect 11152 7148 11204 7200
rect 11428 7148 11480 7200
rect 14740 7284 14792 7336
rect 15200 7284 15252 7336
rect 13360 7216 13412 7268
rect 14372 7148 14424 7200
rect 14740 7148 14792 7200
rect 16396 7284 16448 7336
rect 16856 7284 16908 7336
rect 15200 7148 15252 7200
rect 15568 7148 15620 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 2872 6944 2924 6996
rect 5540 6944 5592 6996
rect 7748 6944 7800 6996
rect 9864 6944 9916 6996
rect 10600 6944 10652 6996
rect 3424 6808 3476 6860
rect 7104 6876 7156 6928
rect 8116 6876 8168 6928
rect 9404 6876 9456 6928
rect 12716 6944 12768 6996
rect 13636 6944 13688 6996
rect 14280 6944 14332 6996
rect 15752 6944 15804 6996
rect 11888 6919 11940 6928
rect 11888 6885 11897 6919
rect 11897 6885 11931 6919
rect 11931 6885 11940 6919
rect 11888 6876 11940 6885
rect 5356 6604 5408 6656
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 6000 6808 6052 6860
rect 6184 6808 6236 6860
rect 10600 6808 10652 6860
rect 11428 6808 11480 6860
rect 11704 6808 11756 6860
rect 11796 6808 11848 6860
rect 15844 6876 15896 6928
rect 16856 6876 16908 6928
rect 7104 6740 7156 6792
rect 6552 6672 6604 6724
rect 6276 6604 6328 6656
rect 6644 6604 6696 6656
rect 6828 6604 6880 6656
rect 7380 6783 7432 6792
rect 7380 6749 7389 6783
rect 7389 6749 7423 6783
rect 7423 6749 7432 6783
rect 7380 6740 7432 6749
rect 7748 6740 7800 6792
rect 8208 6740 8260 6792
rect 10048 6740 10100 6792
rect 10784 6740 10836 6792
rect 11336 6740 11388 6792
rect 11980 6740 12032 6792
rect 13820 6740 13872 6792
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 14924 6740 14976 6792
rect 15108 6783 15160 6792
rect 15108 6749 15117 6783
rect 15117 6749 15151 6783
rect 15151 6749 15160 6783
rect 15108 6740 15160 6749
rect 16212 6808 16264 6860
rect 15292 6783 15344 6792
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 15476 6783 15528 6792
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 8116 6672 8168 6724
rect 10968 6672 11020 6724
rect 16948 6672 17000 6724
rect 17684 6672 17736 6724
rect 7656 6604 7708 6656
rect 12164 6604 12216 6656
rect 13544 6604 13596 6656
rect 14556 6604 14608 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2872 6375 2924 6384
rect 2872 6341 2881 6375
rect 2881 6341 2915 6375
rect 2915 6341 2924 6375
rect 2872 6332 2924 6341
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 3792 6307 3844 6316
rect 3792 6273 3801 6307
rect 3801 6273 3835 6307
rect 3835 6273 3844 6307
rect 3792 6264 3844 6273
rect 6184 6400 6236 6452
rect 6828 6400 6880 6452
rect 7104 6400 7156 6452
rect 8116 6400 8168 6452
rect 10324 6400 10376 6452
rect 11888 6400 11940 6452
rect 12164 6443 12216 6452
rect 12164 6409 12173 6443
rect 12173 6409 12207 6443
rect 12207 6409 12216 6443
rect 12164 6400 12216 6409
rect 12256 6400 12308 6452
rect 5264 6332 5316 6384
rect 4068 6239 4120 6248
rect 4068 6205 4077 6239
rect 4077 6205 4111 6239
rect 4111 6205 4120 6239
rect 4068 6196 4120 6205
rect 3056 6103 3108 6112
rect 3056 6069 3065 6103
rect 3065 6069 3099 6103
rect 3099 6069 3108 6103
rect 3056 6060 3108 6069
rect 3700 6060 3752 6112
rect 3884 6103 3936 6112
rect 3884 6069 3893 6103
rect 3893 6069 3927 6103
rect 3927 6069 3936 6103
rect 3884 6060 3936 6069
rect 5172 6307 5224 6316
rect 5172 6273 5181 6307
rect 5181 6273 5215 6307
rect 5215 6273 5224 6307
rect 5172 6264 5224 6273
rect 5356 6307 5408 6316
rect 5356 6273 5365 6307
rect 5365 6273 5399 6307
rect 5399 6273 5408 6307
rect 5356 6264 5408 6273
rect 5632 6332 5684 6384
rect 5264 6196 5316 6248
rect 6000 6307 6052 6316
rect 6000 6273 6009 6307
rect 6009 6273 6043 6307
rect 6043 6273 6052 6307
rect 6000 6264 6052 6273
rect 6552 6332 6604 6384
rect 7012 6332 7064 6384
rect 7380 6332 7432 6384
rect 7564 6332 7616 6384
rect 6644 6264 6696 6316
rect 5816 6196 5868 6248
rect 6460 6196 6512 6248
rect 7656 6307 7708 6316
rect 7656 6273 7665 6307
rect 7665 6273 7699 6307
rect 7699 6273 7708 6307
rect 7656 6264 7708 6273
rect 7932 6307 7984 6316
rect 7932 6273 7941 6307
rect 7941 6273 7975 6307
rect 7975 6273 7984 6307
rect 7932 6264 7984 6273
rect 8116 6307 8168 6316
rect 8116 6273 8125 6307
rect 8125 6273 8159 6307
rect 8159 6273 8168 6307
rect 8116 6264 8168 6273
rect 8208 6264 8260 6316
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 7656 6128 7708 6180
rect 8484 6196 8536 6248
rect 9128 6307 9180 6316
rect 9128 6273 9137 6307
rect 9137 6273 9171 6307
rect 9171 6273 9180 6307
rect 9128 6264 9180 6273
rect 9404 6307 9456 6316
rect 9404 6273 9413 6307
rect 9413 6273 9447 6307
rect 9447 6273 9456 6307
rect 9404 6264 9456 6273
rect 8116 6128 8168 6180
rect 8944 6128 8996 6180
rect 9312 6196 9364 6248
rect 9864 6307 9916 6316
rect 9864 6273 9873 6307
rect 9873 6273 9907 6307
rect 9907 6273 9916 6307
rect 9864 6264 9916 6273
rect 9588 6196 9640 6248
rect 10416 6264 10468 6316
rect 10600 6307 10652 6316
rect 10600 6273 10609 6307
rect 10609 6273 10643 6307
rect 10643 6273 10652 6307
rect 10600 6264 10652 6273
rect 10784 6307 10836 6316
rect 10784 6273 10793 6307
rect 10793 6273 10827 6307
rect 10827 6273 10836 6307
rect 10784 6264 10836 6273
rect 11428 6264 11480 6316
rect 11152 6196 11204 6248
rect 4896 6103 4948 6112
rect 4896 6069 4905 6103
rect 4905 6069 4939 6103
rect 4939 6069 4948 6103
rect 4896 6060 4948 6069
rect 5816 6103 5868 6112
rect 5816 6069 5825 6103
rect 5825 6069 5859 6103
rect 5859 6069 5868 6103
rect 5816 6060 5868 6069
rect 6000 6103 6052 6112
rect 6000 6069 6009 6103
rect 6009 6069 6043 6103
rect 6043 6069 6052 6103
rect 6000 6060 6052 6069
rect 9128 6060 9180 6112
rect 10232 6128 10284 6180
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 12256 6264 12308 6316
rect 12532 6307 12584 6316
rect 12532 6273 12541 6307
rect 12541 6273 12575 6307
rect 12575 6273 12584 6307
rect 12532 6264 12584 6273
rect 14372 6375 14424 6384
rect 14372 6341 14381 6375
rect 14381 6341 14415 6375
rect 14415 6341 14424 6375
rect 14372 6332 14424 6341
rect 12348 6196 12400 6248
rect 13176 6307 13228 6316
rect 13176 6273 13185 6307
rect 13185 6273 13219 6307
rect 13219 6273 13228 6307
rect 13176 6264 13228 6273
rect 13452 6307 13504 6316
rect 13452 6273 13461 6307
rect 13461 6273 13495 6307
rect 13495 6273 13504 6307
rect 13452 6264 13504 6273
rect 13728 6264 13780 6316
rect 14280 6264 14332 6316
rect 14556 6307 14608 6316
rect 14556 6273 14565 6307
rect 14565 6273 14599 6307
rect 14599 6273 14608 6307
rect 14556 6264 14608 6273
rect 15660 6400 15712 6452
rect 15844 6400 15896 6452
rect 16212 6400 16264 6452
rect 17224 6400 17276 6452
rect 15936 6332 15988 6384
rect 17040 6332 17092 6384
rect 15292 6196 15344 6248
rect 9680 6103 9732 6112
rect 9680 6069 9689 6103
rect 9689 6069 9723 6103
rect 9723 6069 9732 6103
rect 9680 6060 9732 6069
rect 10324 6060 10376 6112
rect 14556 6128 14608 6180
rect 14924 6128 14976 6180
rect 10876 6060 10928 6112
rect 11152 6060 11204 6112
rect 11980 6060 12032 6112
rect 12256 6103 12308 6112
rect 12256 6069 12265 6103
rect 12265 6069 12299 6103
rect 12299 6069 12308 6103
rect 12256 6060 12308 6069
rect 12992 6103 13044 6112
rect 12992 6069 13001 6103
rect 13001 6069 13035 6103
rect 13035 6069 13044 6103
rect 12992 6060 13044 6069
rect 14464 6060 14516 6112
rect 15752 6264 15804 6316
rect 16856 6264 16908 6316
rect 17040 6239 17092 6248
rect 17040 6205 17049 6239
rect 17049 6205 17083 6239
rect 17083 6205 17092 6239
rect 17040 6196 17092 6205
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 2872 5856 2924 5908
rect 3608 5856 3660 5908
rect 3700 5856 3752 5908
rect 4804 5899 4856 5908
rect 4804 5865 4813 5899
rect 4813 5865 4847 5899
rect 4847 5865 4856 5899
rect 4804 5856 4856 5865
rect 4896 5856 4948 5908
rect 5172 5856 5224 5908
rect 5816 5856 5868 5908
rect 3516 5720 3568 5772
rect 4436 5763 4488 5772
rect 4436 5729 4445 5763
rect 4445 5729 4479 5763
rect 4479 5729 4488 5763
rect 4436 5720 4488 5729
rect 5540 5720 5592 5772
rect 6000 5720 6052 5772
rect 2504 5584 2556 5636
rect 3884 5695 3936 5704
rect 3884 5661 3926 5695
rect 3926 5661 3936 5695
rect 3884 5652 3936 5661
rect 4988 5695 5040 5704
rect 4988 5661 4997 5695
rect 4997 5661 5031 5695
rect 5031 5661 5040 5695
rect 4988 5652 5040 5661
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 3056 5516 3108 5568
rect 3700 5516 3752 5568
rect 4620 5584 4672 5636
rect 5172 5584 5224 5636
rect 5724 5695 5776 5704
rect 5724 5661 5733 5695
rect 5733 5661 5767 5695
rect 5767 5661 5776 5695
rect 5724 5652 5776 5661
rect 5908 5695 5960 5704
rect 5908 5661 5917 5695
rect 5917 5661 5951 5695
rect 5951 5661 5960 5695
rect 5908 5652 5960 5661
rect 6460 5720 6512 5772
rect 6828 5720 6880 5772
rect 7748 5788 7800 5840
rect 6644 5652 6696 5704
rect 9312 5856 9364 5908
rect 9404 5856 9456 5908
rect 7104 5695 7156 5704
rect 7104 5661 7113 5695
rect 7113 5661 7147 5695
rect 7147 5661 7156 5695
rect 7104 5652 7156 5661
rect 7564 5652 7616 5704
rect 8208 5695 8260 5704
rect 8208 5661 8217 5695
rect 8217 5661 8251 5695
rect 8251 5661 8260 5695
rect 8208 5652 8260 5661
rect 4988 5516 5040 5568
rect 5356 5516 5408 5568
rect 7380 5584 7432 5636
rect 11612 5856 11664 5908
rect 12348 5856 12400 5908
rect 13176 5856 13228 5908
rect 13268 5899 13320 5908
rect 13268 5865 13277 5899
rect 13277 5865 13311 5899
rect 13311 5865 13320 5899
rect 13268 5856 13320 5865
rect 8484 5652 8536 5704
rect 9680 5720 9732 5772
rect 9036 5652 9088 5704
rect 8760 5584 8812 5636
rect 9496 5695 9548 5704
rect 9496 5661 9505 5695
rect 9505 5661 9539 5695
rect 9539 5661 9548 5695
rect 9496 5652 9548 5661
rect 10232 5720 10284 5772
rect 9864 5516 9916 5568
rect 10048 5652 10100 5704
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 10324 5695 10376 5704
rect 10324 5661 10338 5695
rect 10338 5661 10372 5695
rect 10372 5661 10376 5695
rect 10324 5652 10376 5661
rect 10600 5695 10652 5704
rect 10600 5661 10609 5695
rect 10609 5661 10643 5695
rect 10643 5661 10652 5695
rect 10600 5652 10652 5661
rect 11796 5788 11848 5840
rect 12072 5788 12124 5840
rect 13084 5788 13136 5840
rect 15108 5856 15160 5908
rect 15752 5856 15804 5908
rect 10876 5695 10928 5704
rect 10876 5661 10885 5695
rect 10885 5661 10919 5695
rect 10919 5661 10928 5695
rect 10876 5652 10928 5661
rect 11244 5652 11296 5704
rect 10692 5584 10744 5636
rect 11428 5652 11480 5704
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 11796 5652 11848 5661
rect 11980 5695 12032 5704
rect 11980 5661 11989 5695
rect 11989 5661 12023 5695
rect 12023 5661 12032 5695
rect 11980 5652 12032 5661
rect 11336 5516 11388 5568
rect 12440 5695 12492 5704
rect 12440 5661 12449 5695
rect 12449 5661 12483 5695
rect 12483 5661 12492 5695
rect 12440 5652 12492 5661
rect 13544 5720 13596 5772
rect 13636 5695 13688 5704
rect 13636 5661 13648 5695
rect 13648 5661 13682 5695
rect 13682 5661 13688 5695
rect 13636 5652 13688 5661
rect 14924 5695 14976 5704
rect 14924 5661 14933 5695
rect 14933 5661 14967 5695
rect 14967 5661 14976 5695
rect 14924 5652 14976 5661
rect 15108 5695 15160 5704
rect 15108 5661 15117 5695
rect 15117 5661 15151 5695
rect 15151 5661 15160 5695
rect 15108 5652 15160 5661
rect 15384 5652 15436 5704
rect 16120 5720 16172 5772
rect 16856 5720 16908 5772
rect 17408 5652 17460 5704
rect 14372 5584 14424 5636
rect 12900 5516 12952 5568
rect 13636 5559 13688 5568
rect 13636 5525 13645 5559
rect 13645 5525 13679 5559
rect 13679 5525 13688 5559
rect 13636 5516 13688 5525
rect 13820 5559 13872 5568
rect 13820 5525 13829 5559
rect 13829 5525 13863 5559
rect 13863 5525 13872 5559
rect 13820 5516 13872 5525
rect 15200 5627 15252 5636
rect 15200 5593 15209 5627
rect 15209 5593 15243 5627
rect 15243 5593 15252 5627
rect 15200 5584 15252 5593
rect 16764 5584 16816 5636
rect 15476 5559 15528 5568
rect 15476 5525 15485 5559
rect 15485 5525 15519 5559
rect 15519 5525 15528 5559
rect 15476 5516 15528 5525
rect 16672 5516 16724 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 4068 5312 4120 5364
rect 6828 5312 6880 5364
rect 2044 5244 2096 5296
rect 3792 5176 3844 5228
rect 6644 5176 6696 5228
rect 4804 5108 4856 5160
rect 6920 5219 6972 5228
rect 6920 5185 6929 5219
rect 6929 5185 6963 5219
rect 6963 5185 6972 5219
rect 6920 5176 6972 5185
rect 7564 5244 7616 5296
rect 8208 5312 8260 5364
rect 8760 5312 8812 5364
rect 8944 5244 8996 5296
rect 7104 5219 7156 5228
rect 7104 5185 7113 5219
rect 7113 5185 7147 5219
rect 7147 5185 7156 5219
rect 7104 5176 7156 5185
rect 8576 5176 8628 5228
rect 8852 5219 8904 5228
rect 8852 5185 8861 5219
rect 8861 5185 8895 5219
rect 8895 5185 8904 5219
rect 8852 5176 8904 5185
rect 11060 5244 11112 5296
rect 13820 5312 13872 5364
rect 10416 5176 10468 5228
rect 10692 5176 10744 5228
rect 8668 5108 8720 5160
rect 8760 5151 8812 5160
rect 8760 5117 8769 5151
rect 8769 5117 8803 5151
rect 8803 5117 8812 5151
rect 8760 5108 8812 5117
rect 4436 5040 4488 5092
rect 5448 4972 5500 5024
rect 5632 5040 5684 5092
rect 11336 5108 11388 5160
rect 14556 5312 14608 5364
rect 14188 5287 14240 5296
rect 14188 5253 14197 5287
rect 14197 5253 14231 5287
rect 14231 5253 14240 5287
rect 14188 5244 14240 5253
rect 15476 5244 15528 5296
rect 12256 5176 12308 5228
rect 12532 5219 12584 5228
rect 12532 5185 12541 5219
rect 12541 5185 12575 5219
rect 12575 5185 12584 5219
rect 12532 5176 12584 5185
rect 12716 5219 12768 5228
rect 12716 5185 12725 5219
rect 12725 5185 12759 5219
rect 12759 5185 12768 5219
rect 12716 5176 12768 5185
rect 13084 5176 13136 5228
rect 13544 5176 13596 5228
rect 9864 5040 9916 5092
rect 10784 5040 10836 5092
rect 7012 4972 7064 5024
rect 7288 4972 7340 5024
rect 7380 5015 7432 5024
rect 7380 4981 7389 5015
rect 7389 4981 7423 5015
rect 7423 4981 7432 5015
rect 7380 4972 7432 4981
rect 11244 4972 11296 5024
rect 12348 5015 12400 5024
rect 12348 4981 12357 5015
rect 12357 4981 12391 5015
rect 12391 4981 12400 5015
rect 12348 4972 12400 4981
rect 12440 4972 12492 5024
rect 13636 5151 13688 5160
rect 13636 5117 13645 5151
rect 13645 5117 13679 5151
rect 13679 5117 13688 5151
rect 13636 5108 13688 5117
rect 13728 5151 13780 5160
rect 13728 5117 13737 5151
rect 13737 5117 13771 5151
rect 13771 5117 13780 5151
rect 13728 5108 13780 5117
rect 14280 5219 14332 5228
rect 14280 5185 14289 5219
rect 14289 5185 14323 5219
rect 14323 5185 14332 5219
rect 14280 5176 14332 5185
rect 15292 5219 15344 5228
rect 15292 5185 15301 5219
rect 15301 5185 15335 5219
rect 15335 5185 15344 5219
rect 15292 5176 15344 5185
rect 15752 5312 15804 5364
rect 16028 5244 16080 5296
rect 16672 5312 16724 5364
rect 16212 5219 16264 5228
rect 16212 5185 16221 5219
rect 16221 5185 16255 5219
rect 16255 5185 16264 5219
rect 16212 5176 16264 5185
rect 16304 5108 16356 5160
rect 12992 5015 13044 5024
rect 12992 4981 13001 5015
rect 13001 4981 13035 5015
rect 13035 4981 13044 5015
rect 12992 4972 13044 4981
rect 13912 4972 13964 5024
rect 15200 5040 15252 5092
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 5540 4768 5592 4820
rect 3424 4700 3476 4752
rect 5356 4700 5408 4752
rect 8760 4768 8812 4820
rect 9956 4768 10008 4820
rect 10600 4768 10652 4820
rect 11336 4811 11388 4820
rect 11336 4777 11345 4811
rect 11345 4777 11379 4811
rect 11379 4777 11388 4811
rect 11336 4768 11388 4777
rect 4712 4564 4764 4616
rect 5816 4632 5868 4684
rect 7196 4700 7248 4752
rect 12348 4768 12400 4820
rect 13452 4768 13504 4820
rect 14832 4768 14884 4820
rect 15752 4811 15804 4820
rect 15752 4777 15761 4811
rect 15761 4777 15795 4811
rect 15795 4777 15804 4811
rect 15752 4768 15804 4777
rect 15936 4811 15988 4820
rect 15936 4777 15945 4811
rect 15945 4777 15979 4811
rect 15979 4777 15988 4811
rect 15936 4768 15988 4777
rect 5908 4607 5960 4616
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 3148 4496 3200 4548
rect 5356 4496 5408 4548
rect 6828 4607 6880 4616
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 6920 4607 6972 4616
rect 6920 4573 6929 4607
rect 6929 4573 6963 4607
rect 6963 4573 6972 4607
rect 6920 4564 6972 4573
rect 7012 4564 7064 4616
rect 7380 4607 7432 4616
rect 7380 4573 7389 4607
rect 7389 4573 7423 4607
rect 7423 4573 7432 4607
rect 7380 4564 7432 4573
rect 7472 4607 7524 4616
rect 7472 4573 7481 4607
rect 7481 4573 7515 4607
rect 7515 4573 7524 4607
rect 7472 4564 7524 4573
rect 7840 4564 7892 4616
rect 11428 4675 11480 4684
rect 11428 4641 11437 4675
rect 11437 4641 11471 4675
rect 11471 4641 11480 4675
rect 13268 4700 13320 4752
rect 14464 4700 14516 4752
rect 14740 4700 14792 4752
rect 11428 4632 11480 4641
rect 11520 4607 11572 4616
rect 11520 4573 11529 4607
rect 11529 4573 11563 4607
rect 11563 4573 11572 4607
rect 11520 4564 11572 4573
rect 13636 4632 13688 4684
rect 5632 4428 5684 4480
rect 6644 4428 6696 4480
rect 7104 4428 7156 4480
rect 7380 4428 7432 4480
rect 11336 4496 11388 4548
rect 13268 4607 13320 4616
rect 13268 4573 13277 4607
rect 13277 4573 13311 4607
rect 13311 4573 13320 4607
rect 13268 4564 13320 4573
rect 13452 4607 13504 4616
rect 13452 4573 13461 4607
rect 13461 4573 13495 4607
rect 13495 4573 13504 4607
rect 13452 4564 13504 4573
rect 13820 4607 13872 4616
rect 13820 4573 13829 4607
rect 13829 4573 13863 4607
rect 13863 4573 13872 4607
rect 13820 4564 13872 4573
rect 15660 4675 15712 4684
rect 15660 4641 15669 4675
rect 15669 4641 15703 4675
rect 15703 4641 15712 4675
rect 15660 4632 15712 4641
rect 16304 4607 16356 4616
rect 11796 4539 11848 4548
rect 11796 4505 11805 4539
rect 11805 4505 11839 4539
rect 11839 4505 11848 4539
rect 11796 4496 11848 4505
rect 11980 4471 12032 4480
rect 11980 4437 12005 4471
rect 12005 4437 12032 4471
rect 11980 4428 12032 4437
rect 13360 4471 13412 4480
rect 13360 4437 13369 4471
rect 13369 4437 13403 4471
rect 13403 4437 13412 4471
rect 13360 4428 13412 4437
rect 14096 4496 14148 4548
rect 16304 4573 16313 4607
rect 16313 4573 16347 4607
rect 16347 4573 16356 4607
rect 16304 4564 16356 4573
rect 16120 4496 16172 4548
rect 14188 4471 14240 4480
rect 14188 4437 14197 4471
rect 14197 4437 14231 4471
rect 14231 4437 14240 4471
rect 14188 4428 14240 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 5908 4224 5960 4276
rect 8576 4267 8628 4276
rect 8576 4233 8585 4267
rect 8585 4233 8619 4267
rect 8619 4233 8628 4267
rect 8576 4224 8628 4233
rect 10324 4224 10376 4276
rect 10968 4267 11020 4276
rect 10968 4233 10977 4267
rect 10977 4233 11011 4267
rect 11011 4233 11020 4267
rect 10968 4224 11020 4233
rect 11152 4224 11204 4276
rect 11796 4224 11848 4276
rect 3792 4156 3844 4208
rect 4712 4199 4764 4208
rect 4712 4165 4721 4199
rect 4721 4165 4755 4199
rect 4755 4165 4764 4199
rect 4712 4156 4764 4165
rect 5632 4156 5684 4208
rect 6644 4199 6696 4208
rect 6644 4165 6653 4199
rect 6653 4165 6687 4199
rect 6687 4165 6696 4199
rect 6644 4156 6696 4165
rect 6828 4156 6880 4208
rect 8484 4156 8536 4208
rect 3148 4131 3200 4140
rect 3148 4097 3157 4131
rect 3157 4097 3191 4131
rect 3191 4097 3200 4131
rect 3148 4088 3200 4097
rect 3424 4131 3476 4140
rect 3424 4097 3433 4131
rect 3433 4097 3467 4131
rect 3467 4097 3476 4131
rect 3424 4088 3476 4097
rect 5724 4088 5776 4140
rect 5816 4131 5868 4140
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 7012 4088 7064 4140
rect 5264 4020 5316 4072
rect 7380 4131 7432 4140
rect 7380 4097 7389 4131
rect 7389 4097 7423 4131
rect 7423 4097 7432 4131
rect 7380 4088 7432 4097
rect 8392 4131 8444 4140
rect 8392 4097 8401 4131
rect 8401 4097 8435 4131
rect 8435 4097 8444 4131
rect 8392 4088 8444 4097
rect 7840 4063 7892 4072
rect 7840 4029 7849 4063
rect 7849 4029 7883 4063
rect 7883 4029 7892 4063
rect 7840 4020 7892 4029
rect 6920 3952 6972 4004
rect 5448 3884 5500 3936
rect 6276 3884 6328 3936
rect 6828 3884 6880 3936
rect 8024 4063 8076 4072
rect 8024 4029 8033 4063
rect 8033 4029 8067 4063
rect 8067 4029 8076 4063
rect 8024 4020 8076 4029
rect 8116 4020 8168 4072
rect 8944 4088 8996 4140
rect 9036 3952 9088 4004
rect 9220 4131 9272 4140
rect 9220 4097 9229 4131
rect 9229 4097 9263 4131
rect 9263 4097 9272 4131
rect 9220 4088 9272 4097
rect 9588 4131 9640 4140
rect 9588 4097 9597 4131
rect 9597 4097 9631 4131
rect 9631 4097 9640 4131
rect 9588 4088 9640 4097
rect 9772 4131 9824 4140
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 9772 4088 9824 4097
rect 9864 4131 9916 4140
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 10692 4156 10744 4208
rect 11980 4267 12032 4276
rect 11980 4233 11989 4267
rect 11989 4233 12023 4267
rect 12023 4233 12032 4267
rect 11980 4224 12032 4233
rect 13084 4267 13136 4276
rect 13084 4233 13093 4267
rect 13093 4233 13127 4267
rect 13127 4233 13136 4267
rect 13084 4224 13136 4233
rect 13268 4224 13320 4276
rect 16212 4224 16264 4276
rect 10508 4088 10560 4140
rect 10784 4131 10836 4140
rect 10784 4097 10793 4131
rect 10793 4097 10827 4131
rect 10827 4097 10836 4131
rect 10784 4088 10836 4097
rect 11704 4131 11756 4140
rect 11704 4097 11713 4131
rect 11713 4097 11747 4131
rect 11747 4097 11756 4131
rect 11704 4088 11756 4097
rect 12072 4088 12124 4140
rect 12164 4131 12216 4140
rect 12164 4097 12173 4131
rect 12173 4097 12207 4131
rect 12207 4097 12216 4131
rect 12164 4088 12216 4097
rect 13360 4199 13412 4208
rect 13360 4165 13369 4199
rect 13369 4165 13403 4199
rect 13403 4165 13412 4199
rect 13360 4156 13412 4165
rect 15016 4199 15068 4208
rect 15016 4165 15025 4199
rect 15025 4165 15059 4199
rect 15059 4165 15068 4199
rect 15016 4156 15068 4165
rect 12624 4020 12676 4072
rect 13268 4131 13320 4140
rect 13268 4097 13277 4131
rect 13277 4097 13311 4131
rect 13311 4097 13320 4131
rect 13268 4088 13320 4097
rect 13544 4088 13596 4140
rect 13728 4131 13780 4140
rect 13728 4097 13737 4131
rect 13737 4097 13771 4131
rect 13771 4097 13780 4131
rect 13728 4088 13780 4097
rect 14372 4088 14424 4140
rect 15200 4088 15252 4140
rect 15660 4131 15712 4140
rect 15660 4097 15669 4131
rect 15669 4097 15703 4131
rect 15703 4097 15712 4131
rect 15660 4088 15712 4097
rect 16120 4156 16172 4208
rect 16304 4088 16356 4140
rect 14188 4020 14240 4072
rect 14280 4020 14332 4072
rect 8300 3884 8352 3936
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 8852 3884 8904 3936
rect 10140 3952 10192 4004
rect 10416 3952 10468 4004
rect 14648 3952 14700 4004
rect 9496 3884 9548 3936
rect 11244 3884 11296 3936
rect 16580 3884 16632 3936
rect 16764 3952 16816 4004
rect 16948 3884 17000 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 5816 3680 5868 3732
rect 7748 3680 7800 3732
rect 7840 3680 7892 3732
rect 8760 3680 8812 3732
rect 3148 3612 3200 3664
rect 5264 3544 5316 3596
rect 7104 3612 7156 3664
rect 9036 3612 9088 3664
rect 9220 3612 9272 3664
rect 9864 3680 9916 3732
rect 10784 3680 10836 3732
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 3516 3476 3568 3528
rect 3976 3408 4028 3460
rect 5356 3519 5408 3528
rect 5356 3485 5365 3519
rect 5365 3485 5399 3519
rect 5399 3485 5408 3519
rect 5356 3476 5408 3485
rect 5448 3519 5500 3528
rect 5448 3485 5457 3519
rect 5457 3485 5491 3519
rect 5491 3485 5500 3519
rect 5448 3476 5500 3485
rect 6552 3519 6604 3528
rect 6552 3485 6561 3519
rect 6561 3485 6595 3519
rect 6595 3485 6604 3519
rect 6552 3476 6604 3485
rect 6736 3476 6788 3528
rect 8484 3544 8536 3596
rect 7104 3451 7156 3460
rect 7104 3417 7113 3451
rect 7113 3417 7147 3451
rect 7147 3417 7156 3451
rect 7104 3408 7156 3417
rect 8576 3476 8628 3528
rect 10692 3544 10744 3596
rect 13820 3680 13872 3732
rect 13544 3612 13596 3664
rect 14280 3612 14332 3664
rect 8852 3408 8904 3460
rect 2780 3340 2832 3392
rect 6000 3340 6052 3392
rect 6276 3340 6328 3392
rect 8944 3340 8996 3392
rect 9312 3340 9364 3392
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 9956 3519 10008 3528
rect 9956 3485 9965 3519
rect 9965 3485 9999 3519
rect 9999 3485 10008 3519
rect 9956 3476 10008 3485
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 9772 3408 9824 3460
rect 10876 3519 10928 3528
rect 10876 3485 10885 3519
rect 10885 3485 10919 3519
rect 10919 3485 10928 3519
rect 10876 3476 10928 3485
rect 11152 3519 11204 3528
rect 11152 3485 11161 3519
rect 11161 3485 11195 3519
rect 11195 3485 11204 3519
rect 11152 3476 11204 3485
rect 11244 3519 11296 3528
rect 11244 3485 11253 3519
rect 11253 3485 11287 3519
rect 11287 3485 11296 3519
rect 11244 3476 11296 3485
rect 11520 3519 11572 3528
rect 11520 3485 11529 3519
rect 11529 3485 11563 3519
rect 11563 3485 11572 3519
rect 11520 3476 11572 3485
rect 11796 3519 11848 3528
rect 11796 3485 11805 3519
rect 11805 3485 11839 3519
rect 11839 3485 11848 3519
rect 11796 3476 11848 3485
rect 12072 3519 12124 3528
rect 12072 3485 12081 3519
rect 12081 3485 12115 3519
rect 12115 3485 12124 3519
rect 12072 3476 12124 3485
rect 11060 3408 11112 3460
rect 13084 3519 13136 3528
rect 13084 3485 13093 3519
rect 13093 3485 13127 3519
rect 13127 3485 13136 3519
rect 13084 3476 13136 3485
rect 10232 3340 10284 3392
rect 12532 3383 12584 3392
rect 12532 3349 12541 3383
rect 12541 3349 12575 3383
rect 12575 3349 12584 3383
rect 12532 3340 12584 3349
rect 13452 3476 13504 3528
rect 14372 3476 14424 3528
rect 14556 3476 14608 3528
rect 15660 3544 15712 3596
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 16120 3476 16172 3528
rect 13636 3408 13688 3460
rect 14648 3408 14700 3460
rect 16580 3408 16632 3460
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 5356 3136 5408 3188
rect 4712 3068 4764 3120
rect 7196 3136 7248 3188
rect 8944 3136 8996 3188
rect 6000 2932 6052 2984
rect 8668 3000 8720 3052
rect 6092 2864 6144 2916
rect 6368 2796 6420 2848
rect 8576 2932 8628 2984
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 9588 3000 9640 3052
rect 9680 2932 9732 2984
rect 9772 2975 9824 2984
rect 9772 2941 9781 2975
rect 9781 2941 9815 2975
rect 9815 2941 9824 2975
rect 9772 2932 9824 2941
rect 10140 3136 10192 3188
rect 10876 3179 10928 3188
rect 10876 3145 10885 3179
rect 10885 3145 10919 3179
rect 10919 3145 10928 3179
rect 10876 3136 10928 3145
rect 12072 3136 12124 3188
rect 12532 3136 12584 3188
rect 10600 3068 10652 3120
rect 12716 3111 12768 3120
rect 12716 3077 12725 3111
rect 12725 3077 12759 3111
rect 12759 3077 12768 3111
rect 12716 3068 12768 3077
rect 12900 3111 12952 3120
rect 12900 3077 12909 3111
rect 12909 3077 12943 3111
rect 12943 3077 12952 3111
rect 12900 3068 12952 3077
rect 10232 3043 10284 3052
rect 10232 3009 10241 3043
rect 10241 3009 10275 3043
rect 10275 3009 10284 3043
rect 10232 3000 10284 3009
rect 10324 3043 10376 3052
rect 10324 3009 10333 3043
rect 10333 3009 10367 3043
rect 10367 3009 10376 3043
rect 10324 3000 10376 3009
rect 10416 3000 10468 3052
rect 10692 3043 10744 3052
rect 10692 3009 10701 3043
rect 10701 3009 10735 3043
rect 10735 3009 10744 3043
rect 10692 3000 10744 3009
rect 11612 3000 11664 3052
rect 7104 2864 7156 2916
rect 7656 2864 7708 2916
rect 11888 2864 11940 2916
rect 13452 3136 13504 3188
rect 15384 3136 15436 3188
rect 13544 3043 13596 3052
rect 13544 3009 13553 3043
rect 13553 3009 13587 3043
rect 13587 3009 13596 3043
rect 13544 3000 13596 3009
rect 13268 2975 13320 2984
rect 13268 2941 13277 2975
rect 13277 2941 13311 2975
rect 13311 2941 13320 2975
rect 13268 2932 13320 2941
rect 13912 2864 13964 2916
rect 11612 2796 11664 2848
rect 12992 2796 13044 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 10232 2592 10284 2644
rect 6828 2431 6880 2440
rect 6828 2397 6837 2431
rect 6837 2397 6871 2431
rect 6871 2397 6880 2431
rect 6828 2388 6880 2397
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 9496 2431 9548 2440
rect 9496 2397 9505 2431
rect 9505 2397 9539 2431
rect 9539 2397 9548 2431
rect 9496 2388 9548 2397
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 12992 2388 13044 2440
rect 6460 2252 6512 2304
rect 9036 2252 9088 2304
rect 9680 2252 9732 2304
rect 13544 2252 13596 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 7746 21026 7802 21704
rect 8390 21026 8446 21704
rect 9678 21026 9734 21704
rect 10322 21026 10378 21704
rect 10966 21026 11022 21704
rect 7746 20998 8064 21026
rect 7746 20904 7802 20998
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 8036 18970 8064 20998
rect 8390 20998 8708 21026
rect 8390 20904 8446 20998
rect 8680 18970 8708 20998
rect 9678 20998 9996 21026
rect 9678 20904 9734 20998
rect 9968 18970 9996 20998
rect 10322 20998 10640 21026
rect 10322 20904 10378 20998
rect 10612 18970 10640 20998
rect 10888 20998 11022 21026
rect 10888 18970 10916 20998
rect 10966 20904 11022 20998
rect 12898 21026 12954 21704
rect 12898 20998 13216 21026
rect 12898 20904 12954 20998
rect 13188 18970 13216 20998
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 8668 18964 8720 18970
rect 8668 18906 8720 18912
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 13176 18964 13228 18970
rect 13176 18906 13228 18912
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 7576 18426 7604 18702
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 5724 17808 5776 17814
rect 5724 17750 5776 17756
rect 2044 17672 2096 17678
rect 2044 17614 2096 17620
rect 2056 15026 2084 17614
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 2516 15026 2544 17478
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5736 17338 5764 17750
rect 7944 17610 7972 18226
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 7932 17604 7984 17610
rect 7932 17546 7984 17552
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 3436 16590 3464 17070
rect 3792 16992 3844 16998
rect 3792 16934 3844 16940
rect 3804 16658 3832 16934
rect 4080 16658 4108 17138
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 3792 16652 3844 16658
rect 4068 16652 4120 16658
rect 3792 16594 3844 16600
rect 3988 16612 4068 16640
rect 2596 16584 2648 16590
rect 2596 16526 2648 16532
rect 3424 16584 3476 16590
rect 3424 16526 3476 16532
rect 2608 16114 2636 16526
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 3068 16153 3096 16458
rect 3054 16144 3110 16153
rect 2596 16108 2648 16114
rect 3054 16079 3056 16088
rect 2596 16050 2648 16056
rect 3108 16079 3110 16088
rect 3056 16050 3108 16056
rect 2608 15502 2636 16050
rect 3068 15706 3096 16050
rect 3332 15972 3384 15978
rect 3332 15914 3384 15920
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 2976 15609 3004 15642
rect 3344 15638 3372 15914
rect 3332 15632 3384 15638
rect 2962 15600 3018 15609
rect 3384 15592 3464 15620
rect 3332 15574 3384 15580
rect 2962 15535 3018 15544
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 848 14544 900 14550
rect 846 14512 848 14521
rect 900 14512 902 14521
rect 846 14447 902 14456
rect 1688 14414 1716 14758
rect 1964 14618 1992 14758
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1492 13728 1544 13734
rect 1490 13696 1492 13705
rect 1544 13696 1546 13705
rect 1490 13631 1546 13640
rect 1596 13326 1624 14010
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1688 12986 1716 13874
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 1964 12986 1992 13126
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1688 8974 1716 9318
rect 1780 8974 1808 9454
rect 1676 8968 1728 8974
rect 1030 8936 1086 8945
rect 1676 8910 1728 8916
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1030 8871 1086 8880
rect 1044 8838 1072 8871
rect 1032 8832 1084 8838
rect 1032 8774 1084 8780
rect 1492 5568 1544 5574
rect 1490 5536 1492 5545
rect 1544 5536 1546 5545
rect 1490 5471 1546 5480
rect 2056 5302 2084 12718
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 2148 10674 2176 10950
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2240 9586 2268 14758
rect 2424 14414 2452 14962
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2516 14260 2544 14962
rect 2424 14232 2544 14260
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2332 13394 2360 13670
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2424 12782 2452 14232
rect 2502 13424 2558 13433
rect 2502 13359 2558 13368
rect 2516 13326 2544 13359
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2608 12866 2636 15438
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2700 14074 2728 14554
rect 2884 14482 2912 14962
rect 2964 14952 3016 14958
rect 3240 14952 3292 14958
rect 2964 14894 3016 14900
rect 3238 14920 3240 14929
rect 3292 14920 3294 14929
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2792 13274 2820 13874
rect 2872 13728 2924 13734
rect 2872 13670 2924 13676
rect 2884 13530 2912 13670
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2872 13320 2924 13326
rect 2700 13246 2820 13274
rect 2870 13288 2872 13297
rect 2924 13288 2926 13297
rect 2700 12986 2728 13246
rect 2870 13223 2926 13232
rect 2872 13184 2924 13190
rect 2778 13152 2834 13161
rect 2872 13126 2924 13132
rect 2778 13087 2834 13096
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2608 12838 2728 12866
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2608 11150 2636 11698
rect 2700 11694 2728 12838
rect 2792 12434 2820 13087
rect 2884 12918 2912 13126
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2976 12442 3004 14894
rect 3238 14855 3294 14864
rect 3252 14822 3280 14855
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 3240 14544 3292 14550
rect 3240 14486 3292 14492
rect 3252 14006 3280 14486
rect 3240 14000 3292 14006
rect 3240 13942 3292 13948
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 3068 13394 3096 13874
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 3148 13320 3200 13326
rect 3146 13288 3148 13297
rect 3200 13288 3202 13297
rect 3146 13223 3202 13232
rect 3252 12968 3280 13942
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3344 12986 3372 13466
rect 3160 12940 3280 12968
rect 3332 12980 3384 12986
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 3068 12617 3096 12786
rect 3160 12782 3188 12940
rect 3332 12922 3384 12928
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3054 12608 3110 12617
rect 3054 12543 3110 12552
rect 2964 12436 3016 12442
rect 2792 12406 2912 12434
rect 2884 12322 2912 12406
rect 2964 12378 3016 12384
rect 2884 12294 3096 12322
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2884 11694 2912 12038
rect 2976 11898 3004 12174
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2700 11150 2728 11630
rect 2596 11144 2648 11150
rect 2594 11112 2596 11121
rect 2688 11144 2740 11150
rect 2648 11112 2650 11121
rect 2688 11086 2740 11092
rect 2594 11047 2650 11056
rect 2884 10742 2912 11630
rect 2976 11082 3004 11698
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 3068 10470 3096 12294
rect 3252 12238 3280 12718
rect 3344 12374 3372 12786
rect 3332 12368 3384 12374
rect 3332 12310 3384 12316
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3252 11898 3280 12174
rect 3436 12170 3464 15592
rect 3516 15564 3568 15570
rect 3516 15506 3568 15512
rect 3528 15065 3556 15506
rect 3514 15056 3570 15065
rect 3514 14991 3570 15000
rect 3700 15020 3752 15026
rect 3528 12918 3556 14991
rect 3700 14962 3752 14968
rect 3608 13388 3660 13394
rect 3608 13330 3660 13336
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3424 12164 3476 12170
rect 3424 12106 3476 12112
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3252 10674 3280 11834
rect 3436 11762 3464 12106
rect 3528 12102 3556 12582
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3528 11830 3556 12038
rect 3516 11824 3568 11830
rect 3516 11766 3568 11772
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3436 11150 3464 11698
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3436 10742 3464 11086
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 3424 10736 3476 10742
rect 3424 10678 3476 10684
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2424 9518 2452 10066
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 2516 9586 2544 9862
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2332 9178 2360 9454
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2424 9110 2452 9454
rect 2700 9178 2728 9522
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2412 9104 2464 9110
rect 2412 9046 2464 9052
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2516 5642 2544 8910
rect 2792 8906 2820 10202
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3160 10010 3188 10610
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3344 10062 3372 10406
rect 3528 10282 3556 11018
rect 3620 10470 3648 13330
rect 3712 12714 3740 14962
rect 3804 13326 3832 16594
rect 3988 15026 4016 16612
rect 4068 16594 4120 16600
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4528 15700 4580 15706
rect 4528 15642 4580 15648
rect 4436 15428 4488 15434
rect 4436 15370 4488 15376
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 4264 15026 4292 15302
rect 4448 15162 4476 15370
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 3988 14414 4016 14962
rect 4080 14482 4108 14962
rect 4540 14804 4568 15642
rect 4632 15570 4660 17070
rect 4816 16590 4844 17206
rect 6012 17202 6040 17478
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 5816 17196 5868 17202
rect 6000 17196 6052 17202
rect 5868 17156 5948 17184
rect 5816 17138 5868 17144
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 5552 16658 5580 17002
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 5264 16584 5316 16590
rect 5368 16561 5396 16594
rect 5264 16526 5316 16532
rect 5354 16552 5410 16561
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4632 15473 4660 15506
rect 4618 15464 4674 15473
rect 4724 15434 4752 16526
rect 4816 16232 4844 16526
rect 5000 16454 5028 16526
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5276 16250 5304 16526
rect 5354 16487 5410 16496
rect 5264 16244 5316 16250
rect 4816 16204 5212 16232
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 4816 15502 4844 16050
rect 5184 16046 5212 16204
rect 5264 16186 5316 16192
rect 5368 16182 5396 16487
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5356 16176 5408 16182
rect 5262 16144 5318 16153
rect 5356 16118 5408 16124
rect 5262 16079 5318 16088
rect 5276 16046 5304 16079
rect 5080 16040 5132 16046
rect 5078 16008 5080 16017
rect 5172 16040 5224 16046
rect 5132 16008 5134 16017
rect 5172 15982 5224 15988
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 5078 15943 5134 15952
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 5078 15464 5134 15473
rect 4618 15399 4674 15408
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4620 15360 4672 15366
rect 4672 15308 4752 15314
rect 4620 15302 4752 15308
rect 4632 15286 4752 15302
rect 4540 14776 4660 14804
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 4080 14074 4108 14418
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4448 14074 4476 14350
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4540 13938 4568 14214
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4068 13864 4120 13870
rect 4066 13832 4068 13841
rect 4120 13832 4122 13841
rect 4066 13767 4122 13776
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3700 12708 3752 12714
rect 3700 12650 3752 12656
rect 3804 12646 3832 13262
rect 3896 12850 3924 13466
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3896 12306 3924 12378
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 3896 12170 3924 12242
rect 3884 12164 3936 12170
rect 3884 12106 3936 12112
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3700 11008 3752 11014
rect 3804 10996 3832 11698
rect 3752 10968 3832 10996
rect 3700 10950 3752 10956
rect 3608 10464 3660 10470
rect 3712 10452 3740 10950
rect 3792 10600 3844 10606
rect 3896 10588 3924 12106
rect 3988 11354 4016 13670
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4264 12850 4292 13126
rect 4632 12918 4660 14776
rect 4724 14414 4752 15286
rect 4816 14482 4844 15438
rect 5078 15399 5080 15408
rect 5132 15399 5134 15408
rect 5080 15370 5132 15376
rect 5184 15366 5212 15982
rect 5460 15978 5488 16390
rect 5552 16017 5580 16390
rect 5644 16250 5672 16662
rect 5920 16590 5948 17156
rect 6000 17138 6052 17144
rect 7012 16992 7064 16998
rect 7012 16934 7064 16940
rect 7024 16726 7052 16934
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 5908 16584 5960 16590
rect 5908 16526 5960 16532
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 5632 16244 5684 16250
rect 5632 16186 5684 16192
rect 5816 16176 5868 16182
rect 5816 16118 5868 16124
rect 5538 16008 5594 16017
rect 5448 15972 5500 15978
rect 5594 15966 5672 15994
rect 5538 15943 5594 15952
rect 5448 15914 5500 15920
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 4712 14408 4764 14414
rect 4710 14376 4712 14385
rect 4764 14376 4766 14385
rect 4710 14311 4766 14320
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4172 12730 4200 12786
rect 4080 12702 4200 12730
rect 4080 12434 4108 12702
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4160 12436 4212 12442
rect 4080 12406 4160 12434
rect 4160 12378 4212 12384
rect 4632 12374 4660 12582
rect 4068 12368 4120 12374
rect 4068 12310 4120 12316
rect 4620 12368 4672 12374
rect 4620 12310 4672 12316
rect 4080 11762 4108 12310
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4436 12232 4488 12238
rect 4540 12209 4568 12242
rect 4436 12174 4488 12180
rect 4526 12200 4582 12209
rect 4448 11898 4476 12174
rect 4526 12135 4582 12144
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4632 11762 4660 12106
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 3988 10742 4016 11290
rect 4080 11286 4108 11698
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4080 10742 4108 11222
rect 4264 11014 4292 11222
rect 4632 11150 4660 11698
rect 4724 11354 4752 14214
rect 4816 13870 4844 14418
rect 5276 14414 5304 15846
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5368 15026 5396 15098
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5368 14056 5396 14962
rect 5184 14028 5396 14056
rect 5080 14000 5132 14006
rect 5184 13988 5212 14028
rect 5132 13960 5212 13988
rect 5080 13942 5132 13948
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4894 13560 4950 13569
rect 4894 13495 4896 13504
rect 4948 13495 4950 13504
rect 4896 13466 4948 13472
rect 5184 13308 5212 13960
rect 5460 13716 5488 15914
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5552 15065 5580 15438
rect 5538 15056 5594 15065
rect 5538 14991 5594 15000
rect 5540 14884 5592 14890
rect 5540 14826 5592 14832
rect 5368 13688 5488 13716
rect 5184 13280 5304 13308
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 4908 12753 4936 12786
rect 4894 12744 4950 12753
rect 4894 12679 4950 12688
rect 5092 12481 5120 12786
rect 5078 12472 5134 12481
rect 5078 12407 5134 12416
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 5078 11792 5134 11801
rect 5078 11727 5134 11736
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4816 10792 4844 11086
rect 4908 11082 4936 11494
rect 5092 11082 5120 11727
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4816 10764 5212 10792
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4528 10668 4580 10674
rect 4580 10628 4660 10656
rect 4528 10610 4580 10616
rect 3844 10560 3924 10588
rect 3792 10542 3844 10548
rect 3712 10424 3832 10452
rect 3608 10406 3660 10412
rect 3436 10254 3556 10282
rect 3332 10056 3384 10062
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2884 8974 2912 9522
rect 2976 9450 3004 9998
rect 3068 9722 3096 9998
rect 3160 9982 3280 10010
rect 3332 9998 3384 10004
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 3054 9616 3110 9625
rect 3054 9551 3056 9560
rect 3108 9551 3110 9560
rect 3056 9522 3108 9528
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2976 9081 3004 9114
rect 2962 9072 3018 9081
rect 2962 9007 3018 9016
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2780 8900 2832 8906
rect 2780 8842 2832 8848
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 2778 8800 2834 8809
rect 2778 8735 2834 8744
rect 2504 5636 2556 5642
rect 2504 5578 2556 5584
rect 2044 5296 2096 5302
rect 2044 5238 2096 5244
rect 2792 3505 2820 8735
rect 3068 7818 3096 8842
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3160 8537 3188 8774
rect 3146 8528 3202 8537
rect 3146 8463 3202 8472
rect 3056 7812 3108 7818
rect 3056 7754 3108 7760
rect 3252 7546 3280 9982
rect 3344 9761 3372 9998
rect 3330 9752 3386 9761
rect 3330 9687 3386 9696
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3344 9382 3372 9522
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3436 7970 3464 10254
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3528 9568 3556 10066
rect 3620 9722 3648 10406
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 3712 9654 3740 9862
rect 3700 9648 3752 9654
rect 3700 9590 3752 9596
rect 3608 9580 3660 9586
rect 3528 9540 3608 9568
rect 3608 9522 3660 9528
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3344 7942 3464 7970
rect 3528 7954 3556 9318
rect 3620 8090 3648 9522
rect 3804 9500 3832 10424
rect 3896 10169 3924 10560
rect 4066 10568 4122 10577
rect 4066 10503 4122 10512
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3988 10198 4016 10406
rect 3976 10192 4028 10198
rect 3882 10160 3938 10169
rect 3976 10134 4028 10140
rect 3882 10095 3938 10104
rect 3884 9988 3936 9994
rect 3884 9930 3936 9936
rect 3712 9472 3832 9500
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3516 7948 3568 7954
rect 3344 7886 3372 7942
rect 3516 7890 3568 7896
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3252 7342 3280 7482
rect 3436 7410 3464 7822
rect 3528 7410 3556 7890
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2884 7002 2912 7142
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 2884 5914 2912 6326
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 3068 5681 3096 6054
rect 3054 5672 3110 5681
rect 3054 5607 3110 5616
rect 3068 5574 3096 5607
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3160 4554 3188 7210
rect 3436 6866 3464 7346
rect 3528 7274 3556 7346
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3712 7206 3740 9472
rect 3896 9432 3924 9930
rect 3804 9404 3924 9432
rect 3976 9444 4028 9450
rect 3804 9110 3832 9404
rect 3976 9386 4028 9392
rect 3792 9104 3844 9110
rect 3792 9046 3844 9052
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3804 8809 3832 8910
rect 3790 8800 3846 8809
rect 3790 8735 3846 8744
rect 3790 8528 3846 8537
rect 3790 8463 3846 8472
rect 3804 7290 3832 8463
rect 3896 8242 3924 9046
rect 3988 8378 4016 9386
rect 4080 9160 4108 10503
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4264 10130 4292 10202
rect 4434 10160 4490 10169
rect 4252 10124 4304 10130
rect 4434 10095 4490 10104
rect 4252 10066 4304 10072
rect 4448 10062 4476 10095
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 4264 9654 4292 9930
rect 4632 9722 4660 10628
rect 4724 10130 4752 10678
rect 5184 10674 5212 10764
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5000 10577 5028 10610
rect 5276 10588 5304 13280
rect 5368 12102 5396 13688
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5460 12238 5488 13466
rect 5552 12986 5580 14826
rect 5644 14006 5672 15966
rect 5724 15972 5776 15978
rect 5724 15914 5776 15920
rect 5736 14006 5764 15914
rect 5828 15910 5856 16118
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 5828 15502 5856 15846
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5828 14346 5856 15438
rect 5920 15094 5948 16526
rect 6104 16454 6132 16526
rect 6460 16516 6512 16522
rect 6460 16458 6512 16464
rect 6552 16516 6604 16522
rect 6552 16458 6604 16464
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 6012 15706 6040 16050
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 6104 15586 6132 16390
rect 6366 16144 6422 16153
rect 6366 16079 6422 16088
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6104 15558 6224 15586
rect 6288 15570 6316 15846
rect 6090 15464 6146 15473
rect 6090 15399 6092 15408
rect 6144 15399 6146 15408
rect 6092 15370 6144 15376
rect 5908 15088 5960 15094
rect 5908 15030 5960 15036
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 5816 14340 5868 14346
rect 5816 14282 5868 14288
rect 5632 14000 5684 14006
rect 5724 14000 5776 14006
rect 5632 13942 5684 13948
rect 5722 13968 5724 13977
rect 5776 13968 5778 13977
rect 5722 13903 5778 13912
rect 5724 13728 5776 13734
rect 5828 13716 5856 14282
rect 5776 13688 5856 13716
rect 5724 13670 5776 13676
rect 5722 13288 5778 13297
rect 5722 13223 5778 13232
rect 5816 13252 5868 13258
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5552 12434 5580 12922
rect 5552 12406 5672 12434
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5460 11336 5488 12174
rect 5552 11830 5580 12242
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 5368 11308 5488 11336
rect 5368 10656 5396 11308
rect 5552 11234 5580 11766
rect 5460 11206 5580 11234
rect 5460 10810 5488 11206
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5552 10810 5580 11018
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5448 10668 5500 10674
rect 5368 10628 5448 10656
rect 5448 10610 5500 10616
rect 4986 10568 5042 10577
rect 5276 10560 5396 10588
rect 4986 10503 5042 10512
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4816 10266 4844 10406
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4804 10056 4856 10062
rect 4710 10024 4766 10033
rect 4804 9998 4856 10004
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 5262 10024 5318 10033
rect 4710 9959 4766 9968
rect 4724 9926 4752 9959
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4436 9172 4488 9178
rect 4080 9132 4292 9160
rect 4264 8974 4292 9132
rect 4436 9114 4488 9120
rect 4448 9081 4476 9114
rect 4434 9072 4490 9081
rect 4434 9007 4490 9016
rect 4068 8968 4120 8974
rect 4160 8968 4212 8974
rect 4068 8910 4120 8916
rect 4158 8936 4160 8945
rect 4252 8968 4304 8974
rect 4212 8936 4214 8945
rect 4080 8634 4108 8910
rect 4252 8910 4304 8916
rect 4158 8871 4214 8880
rect 4264 8634 4292 8910
rect 4632 8838 4660 9522
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 3988 8350 4108 8378
rect 3976 8288 4028 8294
rect 3896 8236 3976 8242
rect 3896 8230 4028 8236
rect 3896 8214 4016 8230
rect 3988 7886 4016 8214
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3884 7404 3936 7410
rect 3988 7392 4016 7822
rect 4080 7410 4108 8350
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4344 8016 4396 8022
rect 4632 7970 4660 8434
rect 4344 7958 4396 7964
rect 3936 7364 4016 7392
rect 3884 7346 3936 7352
rect 3804 7262 3924 7290
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 4758 3464 6802
rect 3712 6361 3740 7142
rect 3514 6352 3570 6361
rect 3514 6287 3516 6296
rect 3568 6287 3570 6296
rect 3698 6352 3754 6361
rect 3804 6322 3832 7142
rect 3698 6287 3754 6296
rect 3792 6316 3844 6322
rect 3516 6258 3568 6264
rect 3792 6258 3844 6264
rect 3896 6202 3924 7262
rect 3804 6174 3924 6202
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3712 5914 3740 6054
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3620 5817 3648 5850
rect 3606 5808 3662 5817
rect 3516 5772 3568 5778
rect 3606 5743 3662 5752
rect 3516 5714 3568 5720
rect 3528 5658 3556 5714
rect 3528 5630 3740 5658
rect 3712 5574 3740 5630
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3804 5234 3832 6174
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3896 5710 3924 6054
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3424 4752 3476 4758
rect 3424 4694 3476 4700
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 3160 4146 3188 4490
rect 3436 4146 3464 4694
rect 3804 4214 3832 5170
rect 3792 4208 3844 4214
rect 3792 4150 3844 4156
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3160 3670 3188 4082
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 3436 3516 3464 4082
rect 3516 3528 3568 3534
rect 2778 3496 2834 3505
rect 3436 3488 3516 3516
rect 3516 3470 3568 3476
rect 3988 3466 4016 7364
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4356 7206 4384 7958
rect 4540 7942 4660 7970
rect 4540 7886 4568 7942
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4540 7750 4568 7822
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4080 5370 4108 6190
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4448 5098 4476 5714
rect 4632 5642 4660 7822
rect 4724 7410 4752 9862
rect 4816 9518 4844 9998
rect 4908 9926 4936 9998
rect 5262 9959 5318 9968
rect 5276 9926 5304 9959
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 5262 9688 5318 9697
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4908 8974 4936 9658
rect 5262 9623 5318 9632
rect 5172 9580 5224 9586
rect 5276 9568 5304 9623
rect 5224 9540 5304 9568
rect 5172 9522 5224 9528
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 5000 9382 5028 9454
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5092 9110 5120 9454
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4816 8294 4844 8774
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5170 8528 5226 8537
rect 5170 8463 5172 8472
rect 5224 8463 5226 8472
rect 5172 8434 5224 8440
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4816 7886 4844 8230
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5276 6390 5304 9540
rect 5368 7478 5396 10560
rect 5460 10130 5488 10610
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5460 7886 5488 10066
rect 5644 9994 5672 12406
rect 5736 12374 5764 13223
rect 5816 13194 5868 13200
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 5828 11744 5856 13194
rect 6012 12889 6040 14350
rect 5998 12880 6054 12889
rect 5908 12844 5960 12850
rect 6104 12850 6132 15370
rect 6196 14249 6224 15558
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 6274 15464 6330 15473
rect 6274 15399 6330 15408
rect 6288 14346 6316 15399
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 6182 14240 6238 14249
rect 6182 14175 6238 14184
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 6196 13841 6224 13874
rect 6182 13832 6238 13841
rect 6182 13767 6238 13776
rect 6380 13410 6408 16079
rect 6472 15473 6500 16458
rect 6564 15910 6592 16458
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6736 16176 6788 16182
rect 6736 16118 6788 16124
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6564 15706 6592 15846
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6458 15464 6514 15473
rect 6458 15399 6514 15408
rect 6460 15360 6512 15366
rect 6460 15302 6512 15308
rect 6472 14618 6500 15302
rect 6564 14940 6592 15642
rect 6748 15638 6776 16118
rect 6840 16114 6868 16390
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6736 15632 6788 15638
rect 6736 15574 6788 15580
rect 6840 15094 6868 16050
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 7024 15026 7052 16662
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 7116 15978 7144 16526
rect 7104 15972 7156 15978
rect 7104 15914 7156 15920
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 6564 14912 6684 14940
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6656 14414 6684 14912
rect 6828 14816 6880 14822
rect 6826 14784 6828 14793
rect 6880 14784 6882 14793
rect 6826 14719 6882 14728
rect 7024 14414 7052 14962
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 7012 14408 7064 14414
rect 7012 14350 7064 14356
rect 6460 14272 6512 14278
rect 6460 14214 6512 14220
rect 6472 13530 6500 14214
rect 6564 13870 6592 14350
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6460 13524 6512 13530
rect 6460 13466 6512 13472
rect 6380 13382 6592 13410
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6380 12986 6408 13262
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 5998 12815 6054 12824
rect 6092 12844 6144 12850
rect 5908 12786 5960 12792
rect 6092 12786 6144 12792
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 5920 12374 5948 12786
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 5908 12368 5960 12374
rect 5908 12310 5960 12316
rect 5908 11824 5960 11830
rect 5908 11766 5960 11772
rect 5736 11716 5856 11744
rect 5736 11286 5764 11716
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5736 10198 5764 11222
rect 5920 11150 5948 11766
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 6012 11150 6040 11630
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 6090 11112 6146 11121
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5828 10441 5856 11018
rect 5920 10577 5948 11086
rect 5906 10568 5962 10577
rect 5906 10503 5962 10512
rect 5814 10432 5870 10441
rect 5814 10367 5870 10376
rect 6012 10198 6040 11086
rect 6090 11047 6092 11056
rect 6144 11047 6146 11056
rect 6092 11018 6144 11024
rect 6092 10668 6144 10674
rect 6092 10610 6144 10616
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5552 9382 5580 9862
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5356 7336 5408 7342
rect 5354 7304 5356 7313
rect 5408 7304 5410 7313
rect 5354 7239 5410 7248
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5264 6384 5316 6390
rect 4894 6352 4950 6361
rect 5264 6326 5316 6332
rect 5368 6322 5396 6598
rect 4894 6287 4950 6296
rect 5172 6316 5224 6322
rect 4802 6216 4858 6225
rect 4802 6151 4858 6160
rect 4816 5914 4844 6151
rect 4908 6118 4936 6287
rect 5172 6258 5224 6264
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 5184 5914 5212 6258
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 4908 5556 4936 5850
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 5000 5574 5028 5646
rect 5172 5636 5224 5642
rect 5276 5624 5304 6190
rect 5224 5596 5304 5624
rect 5172 5578 5224 5584
rect 4816 5528 4936 5556
rect 4988 5568 5040 5574
rect 4816 5166 4844 5528
rect 4988 5510 5040 5516
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 4436 5092 4488 5098
rect 4436 5034 4488 5040
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4724 4214 4752 4558
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 2778 3431 2834 3440
rect 3976 3460 4028 3466
rect 2792 3398 2820 3431
rect 3976 3402 4028 3408
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 4724 3126 4752 4150
rect 5276 4078 5304 5596
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5368 4758 5396 5510
rect 5460 5030 5488 7822
rect 5552 7342 5580 8842
rect 5644 8022 5672 9930
rect 5736 9897 5764 10134
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5722 9888 5778 9897
rect 5722 9823 5778 9832
rect 5828 9654 5856 10066
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5906 9616 5962 9625
rect 5906 9551 5908 9560
rect 5960 9551 5962 9560
rect 5908 9522 5960 9528
rect 5814 9480 5870 9489
rect 5814 9415 5870 9424
rect 5828 8566 5856 9415
rect 6012 9110 6040 9862
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5816 8560 5868 8566
rect 6000 8560 6052 8566
rect 5816 8502 5868 8508
rect 5998 8528 6000 8537
rect 6052 8528 6054 8537
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5736 7970 5764 8502
rect 5998 8463 6054 8472
rect 6104 8430 6132 10610
rect 6196 10266 6224 12718
rect 6368 12708 6420 12714
rect 6368 12650 6420 12656
rect 6380 12306 6408 12650
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6472 11898 6500 12786
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6288 10742 6316 11222
rect 6472 11132 6500 11834
rect 6380 11104 6500 11132
rect 6276 10736 6328 10742
rect 6276 10678 6328 10684
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6196 8514 6224 10202
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 6288 8650 6316 10134
rect 6380 8786 6408 11104
rect 6564 11082 6592 13382
rect 6656 12594 6684 14350
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6748 12850 6776 14010
rect 6840 13190 6868 14282
rect 6932 14249 6960 14282
rect 6918 14240 6974 14249
rect 6918 14175 6974 14184
rect 7208 14090 7236 17274
rect 8036 17202 8064 17478
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7484 16590 7512 17070
rect 8128 16794 8156 18158
rect 8208 17808 8260 17814
rect 8208 17750 8260 17756
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 7472 16584 7524 16590
rect 8116 16584 8168 16590
rect 7472 16526 7524 16532
rect 7852 16544 8116 16572
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7300 15434 7328 15982
rect 7288 15428 7340 15434
rect 7288 15370 7340 15376
rect 7392 15162 7420 16526
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7392 14822 7420 14962
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7024 14062 7236 14090
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6932 13841 6960 13874
rect 6918 13832 6974 13841
rect 6918 13767 6974 13776
rect 6932 13394 6960 13767
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 7024 13258 7052 14062
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7116 13530 7144 13874
rect 7194 13560 7250 13569
rect 7104 13524 7156 13530
rect 7194 13495 7196 13504
rect 7104 13466 7156 13472
rect 7248 13495 7250 13504
rect 7196 13466 7248 13472
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6748 12714 6776 12786
rect 6920 12776 6972 12782
rect 6918 12744 6920 12753
rect 7104 12776 7156 12782
rect 6972 12744 6974 12753
rect 6736 12708 6788 12714
rect 7104 12718 7156 12724
rect 6918 12679 6974 12688
rect 6736 12650 6788 12656
rect 6656 12566 6868 12594
rect 6736 12436 6788 12442
rect 6840 12434 6868 12566
rect 7116 12434 7144 12718
rect 6840 12406 7144 12434
rect 6736 12378 6788 12384
rect 6748 12306 6776 12378
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6748 11694 6776 12242
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6656 11150 6684 11562
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6748 11286 6776 11494
rect 6736 11280 6788 11286
rect 6932 11257 6960 11494
rect 6736 11222 6788 11228
rect 6918 11248 6974 11257
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6472 9722 6500 10950
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6458 9616 6514 9625
rect 6458 9551 6460 9560
rect 6512 9551 6514 9560
rect 6460 9522 6512 9528
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6472 8974 6500 9318
rect 6564 8974 6592 9862
rect 6656 9625 6684 11086
rect 6642 9616 6698 9625
rect 6642 9551 6698 9560
rect 6748 9500 6776 11222
rect 6918 11183 6974 11192
rect 6828 11144 6880 11150
rect 6826 11112 6828 11121
rect 6920 11144 6972 11150
rect 6880 11112 6882 11121
rect 6920 11086 6972 11092
rect 6826 11047 6882 11056
rect 6932 10810 6960 11086
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7024 10674 7052 12406
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7208 12238 7236 12310
rect 7300 12238 7328 14758
rect 7484 14362 7512 16526
rect 7852 16250 7880 16544
rect 8116 16526 8168 16532
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7852 15978 7880 16050
rect 7564 15972 7616 15978
rect 7564 15914 7616 15920
rect 7840 15972 7892 15978
rect 7840 15914 7892 15920
rect 7576 15502 7604 15914
rect 7746 15600 7802 15609
rect 7746 15535 7802 15544
rect 7760 15502 7788 15535
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7748 15496 7800 15502
rect 7852 15473 7880 15914
rect 7944 15502 7972 16186
rect 8024 15632 8076 15638
rect 8220 15586 8248 17750
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8024 15574 8076 15580
rect 7932 15496 7984 15502
rect 7748 15438 7800 15444
rect 7838 15464 7894 15473
rect 7576 15026 7604 15438
rect 7932 15438 7984 15444
rect 7838 15399 7894 15408
rect 7944 15162 7972 15438
rect 8036 15434 8064 15574
rect 8128 15558 8248 15586
rect 8024 15428 8076 15434
rect 8024 15370 8076 15376
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 8024 15088 8076 15094
rect 8024 15030 8076 15036
rect 7564 15020 7616 15026
rect 7840 15020 7892 15026
rect 7616 14980 7696 15008
rect 7564 14962 7616 14968
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7576 14482 7604 14758
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7668 14414 7696 14980
rect 7840 14962 7892 14968
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 7852 14822 7880 14962
rect 7840 14816 7892 14822
rect 7840 14758 7892 14764
rect 7852 14498 7880 14758
rect 7944 14618 7972 14962
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7852 14470 7972 14498
rect 7392 14334 7512 14362
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 7392 12322 7420 14334
rect 7656 14000 7708 14006
rect 7484 13948 7656 13954
rect 7484 13942 7708 13948
rect 7484 13926 7696 13942
rect 7484 12434 7512 13926
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7484 12406 7604 12434
rect 7392 12294 7512 12322
rect 7484 12238 7512 12294
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7116 11218 7144 12174
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7208 11898 7236 12038
rect 7392 11898 7420 12174
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 7102 10432 7158 10441
rect 6840 10266 6868 10406
rect 7102 10367 7158 10376
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6840 9722 6868 9930
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6656 9472 6776 9500
rect 6828 9512 6880 9518
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6380 8758 6592 8786
rect 6288 8622 6500 8650
rect 6196 8486 6316 8514
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 5736 7942 5856 7970
rect 5828 7886 5856 7942
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5552 7002 5580 7278
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5644 6390 5672 7142
rect 5724 6792 5776 6798
rect 5722 6760 5724 6769
rect 5776 6760 5778 6769
rect 5722 6695 5778 6704
rect 5632 6384 5684 6390
rect 5632 6326 5684 6332
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5552 4826 5580 5714
rect 5644 5098 5672 6326
rect 5736 5794 5764 6695
rect 5828 6254 5856 7822
rect 5920 7750 5948 8366
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 6000 7880 6052 7886
rect 5998 7848 6000 7857
rect 6052 7848 6054 7857
rect 5998 7783 6054 7792
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6012 7478 6040 7686
rect 6000 7472 6052 7478
rect 6000 7414 6052 7420
rect 5998 7032 6054 7041
rect 5998 6967 6054 6976
rect 6012 6866 6040 6967
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6012 6322 6040 6802
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 5828 5914 5856 6054
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5736 5766 5856 5794
rect 6012 5778 6040 6054
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5354 4584 5410 4593
rect 5354 4519 5356 4528
rect 5408 4519 5410 4528
rect 5356 4490 5408 4496
rect 5644 4486 5672 5034
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5644 4214 5672 4422
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 5736 4146 5764 5646
rect 5828 4842 5856 5766
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5920 5409 5948 5646
rect 5906 5400 5962 5409
rect 5906 5335 5962 5344
rect 5828 4814 6040 4842
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5828 4146 5856 4626
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5920 4282 5948 4558
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5276 3602 5304 4014
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5460 3534 5488 3878
rect 5828 3738 5856 4082
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 5368 3194 5396 3470
rect 6012 3398 6040 4814
rect 6104 3602 6132 7958
rect 6196 6866 6224 8298
rect 6288 7970 6316 8486
rect 6288 7942 6408 7970
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6288 7546 6316 7822
rect 6380 7750 6408 7942
rect 6472 7834 6500 8622
rect 6564 8498 6592 8758
rect 6656 8537 6684 9472
rect 6932 9500 6960 10202
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 7024 9586 7052 9862
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6880 9472 6960 9500
rect 6828 9454 6880 9460
rect 6840 9382 6868 9454
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6932 9160 6960 9472
rect 7012 9444 7064 9450
rect 7116 9432 7144 10367
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7300 10062 7328 10202
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7208 9926 7236 9998
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7064 9404 7144 9432
rect 7012 9386 7064 9392
rect 6932 9132 7052 9160
rect 6918 9072 6974 9081
rect 6918 9007 6974 9016
rect 6932 8974 6960 9007
rect 6920 8968 6972 8974
rect 6748 8916 6920 8922
rect 6748 8910 6972 8916
rect 6748 8894 6960 8910
rect 7024 8906 7052 9132
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 7012 8900 7064 8906
rect 6642 8528 6698 8537
rect 6552 8492 6604 8498
rect 6642 8463 6698 8472
rect 6552 8434 6604 8440
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6564 7993 6592 8026
rect 6550 7984 6606 7993
rect 6656 7954 6684 8366
rect 6550 7919 6606 7928
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6472 7806 6684 7834
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6564 7410 6592 7482
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6366 7032 6422 7041
rect 6366 6967 6422 6976
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6196 6458 6224 6802
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6288 3942 6316 6598
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 6012 2990 6040 3334
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 6104 2922 6132 3538
rect 6288 3398 6316 3878
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6380 2961 6408 6967
rect 6472 6361 6500 7142
rect 6564 6730 6592 7346
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6564 6390 6592 6666
rect 6656 6662 6684 7806
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6552 6384 6604 6390
rect 6458 6352 6514 6361
rect 6552 6326 6604 6332
rect 6458 6287 6514 6296
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6472 5778 6500 6190
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6564 3534 6592 6326
rect 6656 6322 6684 6598
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6656 5234 6684 5646
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6656 4486 6684 5170
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6656 4214 6684 4422
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 6748 3534 6776 8894
rect 7012 8842 7064 8848
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6918 8800 6974 8809
rect 6840 8090 6868 8774
rect 6918 8735 6974 8744
rect 6932 8566 6960 8735
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 7024 8498 7052 8842
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6840 6916 6868 8026
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 7546 6960 7686
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 7024 7410 7052 8434
rect 7116 8430 7144 9046
rect 7104 8424 7156 8430
rect 7208 8401 7236 9862
rect 7300 9586 7328 9862
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7392 9382 7420 11154
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7484 9042 7512 12174
rect 7576 11830 7604 12406
rect 7564 11824 7616 11830
rect 7564 11766 7616 11772
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7576 11354 7604 11630
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7564 9988 7616 9994
rect 7564 9930 7616 9936
rect 7576 9761 7604 9930
rect 7562 9752 7618 9761
rect 7562 9687 7618 9696
rect 7668 9602 7696 13670
rect 7746 12608 7802 12617
rect 7746 12543 7802 12552
rect 7760 12442 7788 12543
rect 7852 12442 7880 13806
rect 7944 13258 7972 14470
rect 8036 14346 8064 15030
rect 8024 14340 8076 14346
rect 8024 14282 8076 14288
rect 8128 13938 8156 15558
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8220 15337 8248 15438
rect 8206 15328 8262 15337
rect 8206 15263 8262 15272
rect 8312 15162 8340 16050
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8208 14884 8260 14890
rect 8208 14826 8260 14832
rect 8220 14793 8248 14826
rect 8206 14784 8262 14793
rect 8206 14719 8262 14728
rect 8208 14544 8260 14550
rect 8208 14486 8260 14492
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8036 13530 8064 13874
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 7932 13252 7984 13258
rect 7932 13194 7984 13200
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7840 12232 7892 12238
rect 7944 12220 7972 13194
rect 7892 12192 7972 12220
rect 8024 12232 8076 12238
rect 7840 12174 7892 12180
rect 8024 12174 8076 12180
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7760 11218 7788 12038
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7748 11076 7800 11082
rect 7852 11064 7880 12174
rect 8036 11762 8064 12174
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 8116 11756 8168 11762
rect 8116 11698 8168 11704
rect 8128 11626 8156 11698
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 8116 11620 8168 11626
rect 8116 11562 8168 11568
rect 7944 11529 7972 11562
rect 7930 11520 7986 11529
rect 7930 11455 7986 11464
rect 8220 11150 8248 14486
rect 8312 14414 8340 15098
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8312 11762 8340 12310
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8298 11656 8354 11665
rect 8298 11591 8300 11600
rect 8352 11591 8354 11600
rect 8300 11562 8352 11568
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 7800 11036 7880 11064
rect 7748 11018 7800 11024
rect 7760 9994 7788 11018
rect 7944 10810 7972 11086
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7748 9988 7800 9994
rect 7748 9930 7800 9936
rect 7944 9722 7972 10202
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 7576 9586 7788 9602
rect 7944 9586 7972 9658
rect 7564 9580 7788 9586
rect 7616 9574 7788 9580
rect 7564 9522 7616 9528
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7668 9178 7696 9454
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7472 9036 7524 9042
rect 7524 8996 7604 9024
rect 7472 8978 7524 8984
rect 7288 8424 7340 8430
rect 7104 8366 7156 8372
rect 7194 8392 7250 8401
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 6840 6888 6960 6916
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6840 6458 6868 6598
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6840 5370 6868 5714
rect 6932 5658 6960 6888
rect 7024 6390 7052 7210
rect 7116 6934 7144 8366
rect 7340 8384 7420 8412
rect 7288 8366 7340 8372
rect 7194 8327 7250 8336
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 7116 6798 7144 6870
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 7116 5710 7144 6394
rect 7104 5704 7156 5710
rect 6932 5630 7052 5658
rect 7104 5646 7156 5652
rect 6918 5536 6974 5545
rect 6918 5471 6974 5480
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6932 5234 6960 5471
rect 6920 5228 6972 5234
rect 7024 5216 7052 5630
rect 7104 5228 7156 5234
rect 7024 5188 7104 5216
rect 6920 5170 6972 5176
rect 7104 5170 7156 5176
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 7024 4622 7052 4966
rect 7208 4758 7236 8327
rect 7286 8256 7342 8265
rect 7286 8191 7342 8200
rect 7300 7886 7328 8191
rect 7392 8090 7420 8384
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7300 7478 7328 7686
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7288 7472 7340 7478
rect 7288 7414 7340 7420
rect 7392 7324 7420 7482
rect 7300 7296 7420 7324
rect 7300 5030 7328 7296
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7392 6390 7420 6734
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 7378 5944 7434 5953
rect 7378 5879 7434 5888
rect 7392 5642 7420 5879
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7196 4752 7248 4758
rect 7196 4694 7248 4700
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6840 4214 6868 4558
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6932 4010 6960 4558
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7024 4049 7052 4082
rect 7010 4040 7066 4049
rect 6920 4004 6972 4010
rect 7010 3975 7066 3984
rect 6920 3946 6972 3952
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6366 2952 6422 2961
rect 6092 2916 6144 2922
rect 6366 2887 6422 2896
rect 6092 2858 6144 2864
rect 6380 2854 6408 2887
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 6840 2446 6868 3878
rect 7116 3670 7144 4422
rect 7104 3664 7156 3670
rect 7104 3606 7156 3612
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7116 2922 7144 3402
rect 7208 3194 7236 4694
rect 7392 4622 7420 4966
rect 7484 4622 7512 8298
rect 7576 8022 7604 8996
rect 7760 8498 7788 9574
rect 7932 9580 7984 9586
rect 7852 9540 7932 9568
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7668 8401 7696 8434
rect 7654 8392 7710 8401
rect 7654 8327 7710 8336
rect 7564 8016 7616 8022
rect 7564 7958 7616 7964
rect 7654 7984 7710 7993
rect 7576 6497 7604 7958
rect 7654 7919 7710 7928
rect 7668 7410 7696 7919
rect 7852 7886 7880 9540
rect 7932 9522 7984 9528
rect 8036 9110 8064 11086
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8312 10742 8340 10950
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8024 9104 8076 9110
rect 8128 9081 8156 9318
rect 8024 9046 8076 9052
rect 8114 9072 8170 9081
rect 8114 9007 8170 9016
rect 8128 8974 8156 9007
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 7932 8900 7984 8906
rect 7932 8842 7984 8848
rect 7944 8498 7972 8842
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7760 7002 7788 7346
rect 7852 7342 7880 7482
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7930 6896 7986 6905
rect 7930 6831 7986 6840
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7562 6488 7618 6497
rect 7562 6423 7618 6432
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 7576 5710 7604 6326
rect 7668 6322 7696 6598
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7576 5302 7604 5646
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7392 4146 7420 4422
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7668 2922 7696 6122
rect 7760 5953 7788 6734
rect 7838 6488 7894 6497
rect 7838 6423 7894 6432
rect 7746 5944 7802 5953
rect 7746 5879 7802 5888
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7760 3738 7788 5782
rect 7852 4622 7880 6423
rect 7944 6322 7972 6831
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 8036 4078 8064 8298
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8128 7970 8156 8230
rect 8220 8090 8248 10610
rect 8298 10568 8354 10577
rect 8298 10503 8354 10512
rect 8312 8401 8340 10503
rect 8404 8498 8432 15302
rect 8496 13802 8524 18702
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 8772 17678 8800 18158
rect 8864 17882 8892 18226
rect 9140 18154 9168 18702
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9128 18148 9180 18154
rect 9128 18090 9180 18096
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 8760 17672 8812 17678
rect 8760 17614 8812 17620
rect 8864 17270 8892 17818
rect 9232 17678 9260 18226
rect 9416 17882 9444 18226
rect 9692 18222 9720 18566
rect 10060 18426 10088 18702
rect 11256 18426 11284 18702
rect 12360 18426 12388 18702
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9692 17762 9720 18022
rect 9784 17882 9812 18226
rect 10060 17882 10088 18226
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10704 17882 10732 18158
rect 11716 18154 11744 18226
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 11704 18148 11756 18154
rect 11704 18090 11756 18096
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 9864 17808 9916 17814
rect 9862 17776 9864 17785
rect 9916 17776 9918 17785
rect 9692 17734 9812 17762
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 9784 17610 9812 17734
rect 9862 17711 9918 17720
rect 10506 17776 10562 17785
rect 10506 17711 10562 17720
rect 10600 17740 10652 17746
rect 10520 17610 10548 17711
rect 10600 17682 10652 17688
rect 9772 17604 9824 17610
rect 9772 17546 9824 17552
rect 10416 17604 10468 17610
rect 10416 17546 10468 17552
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 8852 17264 8904 17270
rect 8852 17206 8904 17212
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8588 16726 8616 17138
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8588 15609 8616 16662
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 8772 16289 8800 16526
rect 8758 16280 8814 16289
rect 8758 16215 8814 16224
rect 8864 16114 8892 16934
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8574 15600 8630 15609
rect 8574 15535 8630 15544
rect 8574 14376 8630 14385
rect 8574 14311 8630 14320
rect 8588 13938 8616 14311
rect 8680 14074 8708 15982
rect 8956 15910 8984 17138
rect 9784 17134 9812 17546
rect 10428 17338 10456 17546
rect 10416 17332 10468 17338
rect 10416 17274 10468 17280
rect 10324 17264 10376 17270
rect 10324 17206 10376 17212
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 10140 17196 10192 17202
rect 10192 17156 10272 17184
rect 10140 17138 10192 17144
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9036 17060 9088 17066
rect 9036 17002 9088 17008
rect 9048 16522 9076 17002
rect 9036 16516 9088 16522
rect 9036 16458 9088 16464
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 8944 15904 8996 15910
rect 8942 15872 8944 15881
rect 8996 15872 8998 15881
rect 8942 15807 8998 15816
rect 8942 15600 8998 15609
rect 9048 15570 9076 16118
rect 9140 15910 9168 16390
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 8942 15535 8998 15544
rect 9036 15564 9088 15570
rect 8760 15496 8812 15502
rect 8760 15438 8812 15444
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 8484 13796 8536 13802
rect 8484 13738 8536 13744
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8588 13326 8616 13738
rect 8576 13320 8628 13326
rect 8574 13288 8576 13297
rect 8628 13288 8630 13297
rect 8574 13223 8630 13232
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8588 12434 8616 13126
rect 8496 12406 8616 12434
rect 8496 12374 8524 12406
rect 8484 12368 8536 12374
rect 8588 12345 8616 12406
rect 8484 12310 8536 12316
rect 8574 12336 8630 12345
rect 8574 12271 8630 12280
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8588 12073 8616 12106
rect 8574 12064 8630 12073
rect 8574 11999 8630 12008
rect 8680 11762 8708 14010
rect 8772 13734 8800 15438
rect 8956 14906 8984 15535
rect 9036 15506 9088 15512
rect 8956 14878 9076 14906
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8864 13938 8892 14350
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8852 13456 8904 13462
rect 8852 13398 8904 13404
rect 8864 13258 8892 13398
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8496 8673 8524 11562
rect 8772 11234 8800 12242
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8680 11206 8800 11234
rect 8680 11150 8708 11206
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8588 10606 8616 11086
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8772 10985 8800 11018
rect 8758 10976 8814 10985
rect 8758 10911 8814 10920
rect 8758 10704 8814 10713
rect 8758 10639 8760 10648
rect 8812 10639 8814 10648
rect 8760 10610 8812 10616
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8588 10198 8616 10542
rect 8668 10464 8720 10470
rect 8666 10432 8668 10441
rect 8720 10432 8722 10441
rect 8666 10367 8722 10376
rect 8576 10192 8628 10198
rect 8576 10134 8628 10140
rect 8772 10062 8800 10610
rect 8864 10470 8892 12174
rect 8956 12073 8984 14758
rect 9048 14346 9076 14878
rect 9140 14618 9168 15846
rect 9232 14929 9260 17070
rect 9876 16794 9904 17138
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9678 16688 9734 16697
rect 9600 16658 9678 16674
rect 9588 16652 9678 16658
rect 9640 16646 9678 16652
rect 9678 16623 9734 16632
rect 9588 16594 9640 16600
rect 9312 16584 9364 16590
rect 9772 16584 9824 16590
rect 9312 16526 9364 16532
rect 9692 16544 9772 16572
rect 9324 16114 9352 16526
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9324 16017 9352 16050
rect 9310 16008 9366 16017
rect 9310 15943 9366 15952
rect 9416 15502 9444 16458
rect 9586 16144 9642 16153
rect 9692 16114 9720 16544
rect 9772 16526 9824 16532
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 9968 16232 9996 16526
rect 10244 16454 10272 17156
rect 10336 16590 10364 17206
rect 10612 17202 10640 17682
rect 10888 17678 10916 18022
rect 11520 17876 11572 17882
rect 11520 17818 11572 17824
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10888 17338 10916 17614
rect 11532 17542 11560 17818
rect 11716 17746 11744 18090
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 9784 16204 9996 16232
rect 9586 16079 9642 16088
rect 9680 16108 9732 16114
rect 9600 16046 9628 16079
rect 9680 16050 9732 16056
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9404 15496 9456 15502
rect 9310 15464 9366 15473
rect 9508 15484 9536 15914
rect 9600 15881 9628 15982
rect 9586 15872 9642 15881
rect 9586 15807 9642 15816
rect 9692 15706 9720 16050
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9784 15586 9812 16204
rect 9862 16144 9918 16153
rect 9862 16079 9918 16088
rect 10140 16108 10192 16114
rect 9876 15706 9904 16079
rect 10140 16050 10192 16056
rect 9954 15872 10010 15881
rect 9954 15807 10010 15816
rect 9968 15706 9996 15807
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9692 15570 9812 15586
rect 9680 15564 9812 15570
rect 9732 15558 9812 15564
rect 9680 15506 9732 15512
rect 9588 15496 9640 15502
rect 9508 15456 9588 15484
rect 9404 15438 9456 15444
rect 9588 15438 9640 15444
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9954 15464 10010 15473
rect 9310 15399 9312 15408
rect 9364 15399 9366 15408
rect 9312 15370 9364 15376
rect 9218 14920 9274 14929
rect 9218 14855 9274 14864
rect 9324 14822 9352 15370
rect 9586 15328 9642 15337
rect 9586 15263 9642 15272
rect 9600 15094 9628 15263
rect 9404 15088 9456 15094
rect 9402 15056 9404 15065
rect 9588 15088 9640 15094
rect 9456 15056 9458 15065
rect 9588 15030 9640 15036
rect 9402 14991 9458 15000
rect 9402 14920 9458 14929
rect 9402 14855 9458 14864
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9036 14340 9088 14346
rect 9036 14282 9088 14288
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 8942 12064 8998 12073
rect 8942 11999 8998 12008
rect 8956 11830 8984 11999
rect 8944 11824 8996 11830
rect 8944 11766 8996 11772
rect 8944 11280 8996 11286
rect 8944 11222 8996 11228
rect 8956 10538 8984 11222
rect 8944 10532 8996 10538
rect 8944 10474 8996 10480
rect 8852 10464 8904 10470
rect 9048 10418 9076 13670
rect 9140 12850 9168 14554
rect 9416 14414 9444 14855
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9404 14408 9456 14414
rect 9508 14385 9536 14554
rect 9404 14350 9456 14356
rect 9494 14376 9550 14385
rect 9494 14311 9550 14320
rect 9600 14113 9628 15030
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9692 14385 9720 14554
rect 9678 14376 9734 14385
rect 9678 14311 9734 14320
rect 9586 14104 9642 14113
rect 9642 14048 9720 14056
rect 9586 14039 9720 14048
rect 9600 14028 9720 14039
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9232 13462 9260 13670
rect 9220 13456 9272 13462
rect 9220 13398 9272 13404
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 9324 13258 9352 13330
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9128 12232 9180 12238
rect 9232 12220 9260 12854
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9180 12192 9260 12220
rect 9128 12174 9180 12180
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9140 11558 9168 12038
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9126 11248 9182 11257
rect 9126 11183 9182 11192
rect 9140 11082 9168 11183
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 9232 10713 9260 12192
rect 9324 11914 9352 12786
rect 9416 12102 9444 13874
rect 9600 13376 9628 13874
rect 9692 13569 9720 14028
rect 9784 13818 9812 15438
rect 9954 15399 10010 15408
rect 10048 15428 10100 15434
rect 9968 15366 9996 15399
rect 10048 15370 10100 15376
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 9876 15094 9904 15302
rect 10060 15162 10088 15370
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 9864 15088 9916 15094
rect 9864 15030 9916 15036
rect 9954 14512 10010 14521
rect 9954 14447 10010 14456
rect 9968 14414 9996 14447
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9876 14074 9904 14350
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9862 13968 9918 13977
rect 9862 13903 9864 13912
rect 9916 13903 9918 13912
rect 9864 13874 9916 13880
rect 9784 13790 9904 13818
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9678 13560 9734 13569
rect 9678 13495 9734 13504
rect 9784 13433 9812 13670
rect 9770 13424 9826 13433
rect 9600 13348 9720 13376
rect 9770 13359 9826 13368
rect 9496 13252 9548 13258
rect 9496 13194 9548 13200
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9508 12481 9536 13194
rect 9600 12918 9628 13194
rect 9692 13190 9720 13348
rect 9784 13190 9812 13359
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9692 12918 9720 13126
rect 9784 13025 9812 13126
rect 9770 13016 9826 13025
rect 9770 12951 9826 12960
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9494 12472 9550 12481
rect 9494 12407 9550 12416
rect 9692 12374 9720 12718
rect 9770 12472 9826 12481
rect 9876 12442 9904 13790
rect 9770 12407 9826 12416
rect 9864 12436 9916 12442
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9784 12152 9812 12407
rect 9864 12378 9916 12384
rect 9692 12124 9812 12152
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9324 11886 9444 11914
rect 9416 11762 9444 11886
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9218 10704 9274 10713
rect 9218 10639 9220 10648
rect 9272 10639 9274 10648
rect 9220 10610 9272 10616
rect 8852 10406 8904 10412
rect 8956 10390 9076 10418
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 8576 10056 8628 10062
rect 8574 10024 8576 10033
rect 8760 10056 8812 10062
rect 8628 10024 8630 10033
rect 8760 9998 8812 10004
rect 8574 9959 8630 9968
rect 8574 9888 8630 9897
rect 8574 9823 8630 9832
rect 8482 8664 8538 8673
rect 8482 8599 8538 8608
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8298 8392 8354 8401
rect 8298 8327 8354 8336
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8496 7970 8524 8502
rect 8588 8498 8616 9823
rect 8956 9674 8984 10390
rect 9128 10192 9180 10198
rect 9128 10134 9180 10140
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 8864 9646 8984 9674
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8680 8498 8708 8774
rect 8864 8498 8892 9646
rect 9048 9450 9076 9998
rect 9036 9444 9088 9450
rect 9036 9386 9088 9392
rect 9048 9110 9076 9386
rect 9036 9104 9088 9110
rect 9036 9046 9088 9052
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 8128 7942 8524 7970
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 8128 6730 8156 6870
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8128 6322 8156 6394
rect 8220 6322 8248 6734
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8116 6180 8168 6186
rect 8116 6122 8168 6128
rect 8128 4078 8156 6122
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8220 5370 8248 5646
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 7852 3738 7880 4014
rect 8312 3942 8340 7822
rect 8404 4146 8432 7942
rect 8588 7857 8616 8434
rect 8574 7848 8630 7857
rect 8630 7806 8708 7834
rect 8574 7783 8630 7792
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8496 5817 8524 6190
rect 8482 5808 8538 5817
rect 8482 5743 8538 5752
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8496 4214 8524 5646
rect 8588 5234 8616 6258
rect 8680 5352 8708 7806
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8772 6225 8800 6258
rect 8758 6216 8814 6225
rect 8758 6151 8814 6160
rect 8772 5642 8800 6151
rect 8760 5636 8812 5642
rect 8760 5578 8812 5584
rect 8864 5409 8892 8434
rect 9048 8401 9076 8434
rect 9034 8392 9090 8401
rect 9034 8327 9090 8336
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9140 7290 9168 10134
rect 9232 8498 9260 10406
rect 9324 9738 9352 11698
rect 9416 11218 9444 11698
rect 9692 11694 9720 12124
rect 9770 12064 9826 12073
rect 9770 11999 9826 12008
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9508 11354 9536 11630
rect 9784 11626 9812 11999
rect 9876 11744 9904 12378
rect 9968 12306 9996 14350
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 10060 13326 10088 13398
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 9876 11716 9996 11744
rect 9862 11656 9918 11665
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9772 11620 9824 11626
rect 9862 11591 9918 11600
rect 9772 11562 9824 11568
rect 9600 11529 9628 11562
rect 9876 11558 9904 11591
rect 9680 11552 9732 11558
rect 9586 11520 9642 11529
rect 9864 11552 9916 11558
rect 9680 11494 9732 11500
rect 9770 11520 9826 11529
rect 9586 11455 9642 11464
rect 9692 11393 9720 11494
rect 9864 11494 9916 11500
rect 9770 11455 9826 11464
rect 9678 11384 9734 11393
rect 9496 11348 9548 11354
rect 9678 11319 9734 11328
rect 9496 11290 9548 11296
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9784 11150 9812 11455
rect 9968 11370 9996 11716
rect 10060 11665 10088 12106
rect 10046 11656 10102 11665
rect 10046 11591 10102 11600
rect 9876 11342 9996 11370
rect 9588 11144 9640 11150
rect 9508 11104 9588 11132
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9416 10674 9444 11018
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9508 10606 9536 11104
rect 9772 11144 9824 11150
rect 9588 11086 9640 11092
rect 9692 11104 9772 11132
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9494 10296 9550 10305
rect 9494 10231 9496 10240
rect 9548 10231 9550 10240
rect 9496 10202 9548 10208
rect 9404 10056 9456 10062
rect 9496 10056 9548 10062
rect 9404 9998 9456 10004
rect 9494 10024 9496 10033
rect 9548 10024 9550 10033
rect 9416 9897 9444 9998
rect 9494 9959 9550 9968
rect 9402 9888 9458 9897
rect 9402 9823 9458 9832
rect 9324 9710 9444 9738
rect 9600 9722 9628 10542
rect 9692 9994 9720 11104
rect 9772 11086 9824 11092
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9218 7984 9274 7993
rect 9218 7919 9274 7928
rect 9232 7886 9260 7919
rect 9324 7886 9352 8910
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 8850 5400 8906 5409
rect 8760 5364 8812 5370
rect 8680 5324 8760 5352
rect 8850 5335 8906 5344
rect 8760 5306 8812 5312
rect 8956 5302 8984 6122
rect 9048 5794 9076 7278
rect 9140 7262 9260 7290
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9140 6118 9168 6258
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9048 5766 9168 5794
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8944 5296 8996 5302
rect 8850 5264 8906 5273
rect 8576 5228 8628 5234
rect 8944 5238 8996 5244
rect 8850 5199 8852 5208
rect 8576 5170 8628 5176
rect 8904 5199 8906 5208
rect 8852 5170 8904 5176
rect 8588 4282 8616 5170
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8484 4208 8536 4214
rect 8484 4150 8536 4156
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 8496 3602 8524 4150
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8588 3534 8616 4218
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8588 2990 8616 3470
rect 8680 3097 8708 5102
rect 8772 4826 8800 5102
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8772 3738 8800 3878
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8864 3466 8892 3878
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 8956 3398 8984 4082
rect 9048 4010 9076 5646
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 9048 3670 9076 3946
rect 9036 3664 9088 3670
rect 9036 3606 9088 3612
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8956 3194 8984 3334
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 8666 3088 8722 3097
rect 8666 3023 8668 3032
rect 8720 3023 8722 3032
rect 8668 2994 8720 3000
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 7656 2916 7708 2922
rect 7656 2858 7708 2864
rect 9140 2446 9168 5766
rect 9232 4146 9260 7262
rect 9416 6934 9444 9710
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9508 8498 9536 9114
rect 9600 8838 9628 9658
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9692 9042 9720 9522
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9784 8514 9812 10406
rect 9876 10198 9904 11342
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9876 8974 9904 9386
rect 9968 8974 9996 11222
rect 10152 11150 10180 16050
rect 10244 15065 10272 16390
rect 10230 15056 10286 15065
rect 10428 15026 10456 16934
rect 10612 16658 10640 17138
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 10874 16688 10930 16697
rect 10600 16652 10652 16658
rect 10874 16623 10930 16632
rect 10600 16594 10652 16600
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10520 16046 10548 16526
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 10704 15094 10732 15370
rect 10796 15366 10824 15914
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10888 15144 10916 16623
rect 11072 16250 11100 17070
rect 11428 17060 11480 17066
rect 11428 17002 11480 17008
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11256 16130 11284 16526
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11164 16102 11284 16130
rect 11336 16108 11388 16114
rect 11072 15910 11100 16050
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 10796 15116 10916 15144
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 10230 14991 10286 15000
rect 10416 15020 10468 15026
rect 10244 13841 10272 14991
rect 10416 14962 10468 14968
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 10414 13968 10470 13977
rect 10414 13903 10470 13912
rect 10230 13832 10286 13841
rect 10230 13767 10286 13776
rect 10428 13569 10456 13903
rect 10414 13560 10470 13569
rect 10414 13495 10470 13504
rect 10428 13326 10456 13495
rect 10520 13433 10548 14418
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10600 14000 10652 14006
rect 10600 13942 10652 13948
rect 10506 13424 10562 13433
rect 10506 13359 10562 13368
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10612 12918 10640 13942
rect 10704 13734 10732 14214
rect 10796 13938 10824 15116
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10704 13530 10732 13670
rect 10888 13530 10916 14962
rect 10980 14550 11008 15030
rect 10968 14544 11020 14550
rect 10968 14486 11020 14492
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10968 13456 11020 13462
rect 10968 13398 11020 13404
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10600 12912 10652 12918
rect 10600 12854 10652 12860
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 10244 11529 10272 12242
rect 10336 11762 10364 12378
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10428 11558 10456 12854
rect 10704 12753 10732 13262
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10690 12744 10746 12753
rect 10690 12679 10746 12688
rect 10704 12646 10732 12679
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10796 12481 10824 12786
rect 10782 12472 10838 12481
rect 10980 12434 11008 13398
rect 11072 12646 11100 15846
rect 11164 14414 11192 16102
rect 11336 16050 11388 16056
rect 11348 15745 11376 16050
rect 11334 15736 11390 15745
rect 11334 15671 11390 15680
rect 11440 15042 11468 17002
rect 11348 15014 11468 15042
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 11348 14249 11376 15014
rect 11428 14952 11480 14958
rect 11428 14894 11480 14900
rect 11440 14482 11468 14894
rect 11532 14618 11560 17478
rect 11624 17202 11652 17614
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11624 15910 11652 17138
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11624 15026 11652 15846
rect 11716 15706 11744 17682
rect 11808 17338 11836 18158
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12176 17814 12204 18022
rect 12360 17882 12388 18158
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12164 17808 12216 17814
rect 12164 17750 12216 17756
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11808 17202 11836 17274
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11796 17060 11848 17066
rect 11796 17002 11848 17008
rect 11808 16726 11836 17002
rect 11796 16720 11848 16726
rect 11796 16662 11848 16668
rect 11704 15700 11756 15706
rect 11756 15660 11836 15688
rect 11704 15642 11756 15648
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 11520 14340 11572 14346
rect 11520 14282 11572 14288
rect 11334 14240 11390 14249
rect 11334 14175 11390 14184
rect 11440 14074 11468 14282
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 10782 12407 10838 12416
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10520 11898 10548 12174
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10416 11552 10468 11558
rect 10230 11520 10286 11529
rect 10416 11494 10468 11500
rect 10230 11455 10286 11464
rect 10322 11384 10378 11393
rect 10428 11354 10456 11494
rect 10506 11384 10562 11393
rect 10322 11319 10378 11328
rect 10416 11348 10468 11354
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10060 10674 10088 10746
rect 10152 10713 10180 11086
rect 10138 10704 10194 10713
rect 10048 10668 10100 10674
rect 10138 10639 10194 10648
rect 10232 10668 10284 10674
rect 10048 10610 10100 10616
rect 10232 10610 10284 10616
rect 10060 10520 10088 10610
rect 10140 10532 10192 10538
rect 10060 10492 10140 10520
rect 10060 10130 10088 10492
rect 10140 10474 10192 10480
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 10244 10010 10272 10610
rect 10060 9982 10272 10010
rect 10060 9586 10088 9982
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10048 9580 10100 9586
rect 10100 9540 10180 9568
rect 10048 9522 10100 9528
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9968 8566 9996 8910
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9600 8486 9812 8514
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 9600 8362 9628 8486
rect 9954 8392 10010 8401
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9772 8356 9824 8362
rect 9954 8327 10010 8336
rect 9772 8298 9824 8304
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9508 8022 9536 8230
rect 9496 8016 9548 8022
rect 9496 7958 9548 7964
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7410 9536 7686
rect 9600 7478 9628 7958
rect 9692 7954 9720 8298
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9692 7546 9720 7686
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9404 6928 9456 6934
rect 9404 6870 9456 6876
rect 9416 6474 9444 6870
rect 9324 6446 9444 6474
rect 9324 6254 9352 6446
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9324 5914 9352 6190
rect 9416 5914 9444 6258
rect 9588 6248 9640 6254
rect 9586 6216 9588 6225
rect 9640 6216 9642 6225
rect 9586 6151 9642 6160
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9692 5778 9720 6054
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9508 5409 9536 5646
rect 9494 5400 9550 5409
rect 9494 5335 9550 5344
rect 9784 4298 9812 8298
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9876 7546 9904 7822
rect 9968 7818 9996 8327
rect 10060 7886 10088 9318
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 9956 7812 10008 7818
rect 9956 7754 10008 7760
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9876 6322 9904 6938
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9876 5098 9904 5510
rect 9864 5092 9916 5098
rect 9864 5034 9916 5040
rect 9968 4826 9996 7754
rect 10046 7440 10102 7449
rect 10046 7375 10102 7384
rect 10060 7342 10088 7375
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10060 5710 10088 6734
rect 10152 5710 10180 9540
rect 10244 8498 10272 9862
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10230 8256 10286 8265
rect 10230 8191 10286 8200
rect 10244 7886 10272 8191
rect 10336 7886 10364 11319
rect 10612 11370 10640 12310
rect 10796 12170 10824 12407
rect 10888 12406 11008 12434
rect 10888 12306 10916 12406
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10784 12164 10836 12170
rect 10784 12106 10836 12112
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10562 11342 10640 11370
rect 10506 11319 10562 11328
rect 10416 11290 10468 11296
rect 10520 11014 10548 11319
rect 10704 11218 10732 11494
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10600 10736 10652 10742
rect 10600 10678 10652 10684
rect 10612 10266 10640 10678
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10704 10470 10732 10542
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10598 9752 10654 9761
rect 10598 9687 10654 9696
rect 10414 9344 10470 9353
rect 10414 9279 10470 9288
rect 10428 8974 10456 9279
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10244 6186 10272 7346
rect 10336 7313 10364 7346
rect 10322 7304 10378 7313
rect 10322 7239 10378 7248
rect 10428 6474 10456 8434
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10520 8090 10548 8298
rect 10612 8090 10640 9687
rect 10704 8974 10732 10406
rect 10796 10044 10824 12106
rect 10888 11150 10916 12242
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11072 11937 11100 12174
rect 11058 11928 11114 11937
rect 11164 11914 11192 13466
rect 11348 13161 11376 14010
rect 11532 13734 11560 14282
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11532 13161 11560 13670
rect 11334 13152 11390 13161
rect 11334 13087 11390 13096
rect 11518 13152 11574 13161
rect 11518 13087 11574 13096
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11242 12472 11298 12481
rect 11242 12407 11298 12416
rect 11256 12238 11284 12407
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11256 12102 11284 12174
rect 11348 12152 11376 12650
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11440 12306 11468 12582
rect 11532 12442 11560 12718
rect 11624 12617 11652 12786
rect 11610 12608 11666 12617
rect 11610 12543 11666 12552
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11428 12164 11480 12170
rect 11348 12124 11428 12152
rect 11428 12106 11480 12112
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11164 11886 11284 11914
rect 11058 11863 11114 11872
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 11152 11144 11204 11150
rect 11256 11132 11284 11886
rect 11440 11354 11468 12106
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 11532 11626 11560 12038
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 11428 11144 11480 11150
rect 11256 11104 11428 11132
rect 11152 11086 11204 11092
rect 11428 11086 11480 11092
rect 10888 10810 10916 11086
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10888 10674 10916 10746
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10876 10192 10928 10198
rect 10874 10160 10876 10169
rect 10928 10160 10930 10169
rect 10874 10095 10930 10104
rect 10796 10016 10916 10044
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10704 8294 10732 8434
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10336 6458 10456 6474
rect 10324 6452 10456 6458
rect 10376 6446 10456 6452
rect 10324 6394 10376 6400
rect 10414 6352 10470 6361
rect 10414 6287 10416 6296
rect 10468 6287 10470 6296
rect 10416 6258 10468 6264
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 10324 6112 10376 6118
rect 10244 6060 10324 6066
rect 10244 6054 10376 6060
rect 10244 6038 10364 6054
rect 10244 5778 10272 6038
rect 10322 5808 10378 5817
rect 10232 5772 10284 5778
rect 10322 5743 10378 5752
rect 10232 5714 10284 5720
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9692 4270 9812 4298
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9232 3670 9260 4082
rect 9496 3936 9548 3942
rect 9600 3913 9628 4082
rect 9496 3878 9548 3884
rect 9586 3904 9642 3913
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9324 3058 9352 3334
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9508 2446 9536 3878
rect 9586 3839 9642 3848
rect 9600 3058 9628 3839
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9692 2990 9720 4270
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9784 3466 9812 4082
rect 9876 3738 9904 4082
rect 10152 4010 10180 5646
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 10152 3618 10180 3946
rect 9876 3590 10180 3618
rect 9876 3534 9904 3590
rect 10244 3534 10272 5714
rect 10336 5710 10364 5743
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10336 4282 10364 5646
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10428 4010 10456 5170
rect 10520 4146 10548 7890
rect 10612 7002 10640 8026
rect 10690 7576 10746 7585
rect 10690 7511 10746 7520
rect 10704 7342 10732 7511
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10612 6322 10640 6802
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10612 5545 10640 5646
rect 10704 5642 10732 7278
rect 10796 6798 10824 9454
rect 10888 9042 10916 10016
rect 10980 9586 11008 10950
rect 11058 10704 11114 10713
rect 11164 10674 11192 11086
rect 11058 10639 11114 10648
rect 11152 10668 11204 10674
rect 11072 10470 11100 10639
rect 11152 10610 11204 10616
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11164 10305 11192 10610
rect 11334 10432 11390 10441
rect 11334 10367 11390 10376
rect 11150 10296 11206 10305
rect 11150 10231 11206 10240
rect 11348 10062 11376 10367
rect 11060 10056 11112 10062
rect 11336 10056 11388 10062
rect 11112 10016 11284 10044
rect 11060 9998 11112 10004
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10874 8664 10930 8673
rect 10874 8599 10930 8608
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10888 6610 10916 8599
rect 11072 8498 11100 9318
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11164 8498 11192 8774
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10980 7410 11008 7686
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10966 7168 11022 7177
rect 10966 7103 11022 7112
rect 10980 6730 11008 7103
rect 11072 7018 11100 8434
rect 11256 8378 11284 10016
rect 11336 9998 11388 10004
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11348 8634 11376 8910
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11164 8350 11284 8378
rect 11164 7342 11192 8350
rect 11348 7886 11376 8434
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11256 7546 11284 7822
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11164 7206 11192 7278
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11256 7018 11284 7346
rect 11440 7290 11468 11086
rect 11532 10742 11560 11222
rect 11520 10736 11572 10742
rect 11520 10678 11572 10684
rect 11518 10432 11574 10441
rect 11518 10367 11574 10376
rect 11532 10130 11560 10367
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11532 9722 11560 10066
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11532 9081 11560 9658
rect 11624 9382 11652 12543
rect 11716 12345 11744 13874
rect 11702 12336 11758 12345
rect 11702 12271 11758 12280
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11716 10062 11744 12174
rect 11808 11914 11836 15660
rect 11992 15162 12020 17614
rect 13004 17610 13032 18226
rect 13372 17746 13400 18566
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13556 17814 13584 18226
rect 13544 17808 13596 17814
rect 13544 17750 13596 17756
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 12992 17604 13044 17610
rect 12992 17546 13044 17552
rect 13360 17604 13412 17610
rect 13360 17546 13412 17552
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12070 16688 12126 16697
rect 12268 16658 12296 17138
rect 12070 16623 12126 16632
rect 12256 16652 12308 16658
rect 12084 16182 12112 16623
rect 12256 16594 12308 16600
rect 12268 16182 12296 16594
rect 12452 16522 12480 17274
rect 13372 17202 13400 17546
rect 13648 17338 13676 18226
rect 13728 18148 13780 18154
rect 13728 18090 13780 18096
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13740 17202 13768 18090
rect 14476 18086 14504 18702
rect 14740 18692 14792 18698
rect 14740 18634 14792 18640
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 13832 17746 13860 18022
rect 14188 17808 14240 17814
rect 14188 17750 14240 17756
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 14200 17338 14228 17750
rect 14476 17678 14504 18022
rect 14752 17882 14780 18634
rect 16488 18352 16540 18358
rect 16488 18294 16540 18300
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 14740 17876 14792 17882
rect 14740 17818 14792 17824
rect 15856 17678 15884 18022
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13176 17060 13228 17066
rect 13176 17002 13228 17008
rect 13188 16590 13216 17002
rect 13372 16998 13400 17138
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 12900 16584 12952 16590
rect 12900 16526 12952 16532
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12452 16182 12480 16458
rect 12622 16280 12678 16289
rect 12622 16215 12678 16224
rect 12072 16176 12124 16182
rect 12072 16118 12124 16124
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12440 16176 12492 16182
rect 12440 16118 12492 16124
rect 12532 16176 12584 16182
rect 12532 16118 12584 16124
rect 12164 16108 12216 16114
rect 12164 16050 12216 16056
rect 12176 15366 12204 16050
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 12268 15094 12296 16118
rect 12452 15434 12480 16118
rect 12440 15428 12492 15434
rect 12440 15370 12492 15376
rect 12544 15314 12572 16118
rect 12636 15502 12664 16215
rect 12912 16153 12940 16526
rect 13096 16182 13124 16526
rect 13464 16454 13492 17070
rect 13648 16590 13676 17070
rect 13740 16794 13768 17138
rect 14476 17134 14504 17614
rect 16028 17604 16080 17610
rect 16028 17546 16080 17552
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13740 16674 13768 16730
rect 13740 16646 13860 16674
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13648 16182 13676 16526
rect 13740 16454 13768 16526
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13084 16176 13136 16182
rect 12898 16144 12954 16153
rect 13084 16118 13136 16124
rect 13636 16176 13688 16182
rect 13636 16118 13688 16124
rect 13740 16114 13768 16390
rect 13832 16114 13860 16646
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13924 16454 13952 16594
rect 13912 16448 13964 16454
rect 13912 16390 13964 16396
rect 14108 16114 14136 17070
rect 14648 17060 14700 17066
rect 14648 17002 14700 17008
rect 14280 16244 14332 16250
rect 14280 16186 14332 16192
rect 12898 16079 12954 16088
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 14096 16108 14148 16114
rect 14096 16050 14148 16056
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12452 15286 12572 15314
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 12346 14512 12402 14521
rect 12346 14447 12402 14456
rect 12360 14414 12388 14447
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11886 12880 11942 12889
rect 11992 12850 12020 13738
rect 11886 12815 11888 12824
rect 11940 12815 11942 12824
rect 11980 12844 12032 12850
rect 11888 12786 11940 12792
rect 11980 12786 12032 12792
rect 12176 12186 12204 13806
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12268 12866 12296 13194
rect 12346 13016 12402 13025
rect 12346 12951 12348 12960
rect 12400 12951 12402 12960
rect 12348 12922 12400 12928
rect 12268 12838 12388 12866
rect 12256 12776 12308 12782
rect 12256 12718 12308 12724
rect 11992 12158 12204 12186
rect 11808 11886 11928 11914
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11808 11354 11836 11766
rect 11900 11354 11928 11886
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11992 11234 12020 12158
rect 12268 11937 12296 12718
rect 12360 12714 12388 12838
rect 12348 12708 12400 12714
rect 12348 12650 12400 12656
rect 12360 12238 12388 12650
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12360 12102 12388 12174
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12254 11928 12310 11937
rect 12254 11863 12310 11872
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 11808 11206 12020 11234
rect 11808 10577 11836 11206
rect 11980 11144 12032 11150
rect 12084 11121 12112 11698
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 11980 11086 12032 11092
rect 12070 11112 12126 11121
rect 11886 10840 11942 10849
rect 11992 10810 12020 11086
rect 12070 11047 12126 11056
rect 12176 10996 12204 11562
rect 12268 11558 12296 11863
rect 12348 11688 12400 11694
rect 12452 11665 12480 15286
rect 12808 15088 12860 15094
rect 12806 15056 12808 15065
rect 12860 15056 12862 15065
rect 12532 15020 12584 15026
rect 12806 14991 12862 15000
rect 12532 14962 12584 14968
rect 12544 14618 12572 14962
rect 13096 14958 13124 15982
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13464 15609 13492 15914
rect 13450 15600 13506 15609
rect 13450 15535 13506 15544
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13188 15026 13216 15302
rect 13464 15026 13492 15535
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12728 14482 12756 14758
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12820 14414 12848 14894
rect 12912 14550 12940 14894
rect 13004 14618 13032 14894
rect 12992 14612 13044 14618
rect 12992 14554 13044 14560
rect 12900 14544 12952 14550
rect 12900 14486 12952 14492
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12544 12434 12572 14350
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12728 13190 12756 13670
rect 12912 13462 12940 14282
rect 13096 13938 13124 14894
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 12900 13456 12952 13462
rect 12900 13398 12952 13404
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 12992 13320 13044 13326
rect 12990 13288 12992 13297
rect 13044 13288 13046 13297
rect 12990 13223 13046 13232
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12544 12406 12664 12434
rect 12530 12200 12586 12209
rect 12530 12135 12586 12144
rect 12348 11630 12400 11636
rect 12438 11656 12494 11665
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12360 11218 12388 11630
rect 12544 11626 12572 12135
rect 12438 11591 12494 11600
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12176 10968 12388 10996
rect 11886 10775 11942 10784
rect 11980 10804 12032 10810
rect 11794 10568 11850 10577
rect 11794 10503 11850 10512
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11716 9674 11744 9998
rect 11808 9994 11836 10406
rect 11900 10062 11928 10775
rect 11980 10746 12032 10752
rect 12164 10736 12216 10742
rect 12084 10684 12164 10690
rect 12084 10678 12216 10684
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 12084 10662 12204 10678
rect 11992 10062 12020 10610
rect 12084 10606 12112 10662
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11900 9761 11928 9998
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 11886 9752 11942 9761
rect 11886 9687 11942 9696
rect 11980 9716 12032 9722
rect 11716 9646 11836 9674
rect 11980 9658 12032 9664
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11518 9072 11574 9081
rect 11518 9007 11574 9016
rect 11520 8016 11572 8022
rect 11518 7984 11520 7993
rect 11572 7984 11574 7993
rect 11518 7919 11574 7928
rect 11532 7886 11560 7919
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11520 7472 11572 7478
rect 11520 7414 11572 7420
rect 11532 7313 11560 7414
rect 11072 6990 11284 7018
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10888 6582 11008 6610
rect 10782 6488 10838 6497
rect 10782 6423 10838 6432
rect 10796 6322 10824 6423
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10692 5636 10744 5642
rect 10692 5578 10744 5584
rect 10598 5536 10654 5545
rect 10598 5471 10654 5480
rect 10612 4826 10640 5471
rect 10704 5234 10732 5578
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10704 4214 10732 5170
rect 10796 5098 10824 6258
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10888 5710 10916 6054
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10784 5092 10836 5098
rect 10784 5034 10836 5040
rect 10980 4282 11008 6582
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11164 6118 11192 6190
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11256 5710 11284 6990
rect 11348 7262 11468 7290
rect 11518 7304 11574 7313
rect 11348 6798 11376 7262
rect 11518 7239 11574 7248
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11440 6866 11468 7142
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11348 6361 11376 6734
rect 11334 6352 11390 6361
rect 11334 6287 11390 6296
rect 11428 6316 11480 6322
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11348 5574 11376 6287
rect 11428 6258 11480 6264
rect 11440 5710 11468 6258
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 10692 4208 10744 4214
rect 10598 4176 10654 4185
rect 10508 4140 10560 4146
rect 10692 4150 10744 4156
rect 10598 4111 10654 4120
rect 10508 4082 10560 4088
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 9864 3528 9916 3534
rect 9956 3528 10008 3534
rect 9864 3470 9916 3476
rect 9954 3496 9956 3505
rect 10140 3528 10192 3534
rect 10008 3496 10010 3505
rect 9772 3460 9824 3466
rect 10140 3470 10192 3476
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 9954 3431 10010 3440
rect 9772 3402 9824 3408
rect 10152 3194 10180 3470
rect 10244 3398 10272 3470
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10428 3058 10456 3946
rect 10612 3126 10640 4111
rect 10704 3602 10732 4150
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 10796 3738 10824 4082
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10876 3528 10928 3534
rect 10690 3496 10746 3505
rect 10876 3470 10928 3476
rect 10690 3431 10746 3440
rect 10600 3120 10652 3126
rect 10600 3062 10652 3068
rect 10704 3058 10732 3431
rect 10888 3194 10916 3470
rect 11072 3466 11100 5238
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11164 3534 11192 4218
rect 11256 3942 11284 4966
rect 11348 4826 11376 5102
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11348 4554 11376 4762
rect 11440 4690 11468 5646
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11532 4622 11560 7239
rect 11624 5914 11652 9114
rect 11716 8906 11744 9454
rect 11808 9382 11836 9646
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11796 9104 11848 9110
rect 11796 9046 11848 9052
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11808 8548 11836 9046
rect 11886 8664 11942 8673
rect 11886 8599 11942 8608
rect 11716 8520 11836 8548
rect 11716 7528 11744 8520
rect 11900 8498 11928 8599
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11992 7886 12020 9658
rect 12084 9586 12112 9930
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12084 8106 12112 9318
rect 12176 8294 12204 9930
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12268 9353 12296 9522
rect 12254 9344 12310 9353
rect 12254 9279 12310 9288
rect 12254 9072 12310 9081
rect 12254 9007 12310 9016
rect 12268 8974 12296 9007
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12268 8566 12296 8910
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12084 8078 12204 8106
rect 12072 8016 12124 8022
rect 12072 7958 12124 7964
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11716 7500 11928 7528
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11808 6866 11836 7346
rect 11900 6934 11928 7500
rect 11992 7410 12020 7822
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11888 6928 11940 6934
rect 12084 6905 12112 7958
rect 12176 7954 12204 8078
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12268 7546 12296 7822
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 11888 6870 11940 6876
rect 12070 6896 12126 6905
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11716 6322 11744 6802
rect 11794 6760 11850 6769
rect 11794 6695 11850 6704
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11808 5930 11836 6695
rect 11900 6458 11928 6870
rect 12070 6831 12126 6840
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11716 5902 11836 5930
rect 11716 5760 11744 5902
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11624 5732 11744 5760
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11256 3534 11284 3878
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11520 3528 11572 3534
rect 11624 3516 11652 5732
rect 11808 5710 11836 5782
rect 11796 5704 11848 5710
rect 11716 5664 11796 5692
rect 11716 4146 11744 5664
rect 11796 5646 11848 5652
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11808 4282 11836 4490
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11808 3534 11836 4218
rect 11572 3488 11652 3516
rect 11520 3470 11572 3476
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 11624 3058 11652 3488
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9692 2446 9720 2926
rect 9784 2446 9812 2926
rect 10244 2650 10272 2994
rect 10336 2961 10364 2994
rect 10322 2952 10378 2961
rect 10322 2887 10378 2896
rect 11624 2854 11652 2994
rect 11900 2922 11928 6258
rect 11992 6118 12020 6734
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6458 12204 6598
rect 12268 6458 12296 7346
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12268 6322 12296 6394
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12360 6254 12388 10968
rect 12452 10169 12480 11086
rect 12636 11014 12664 12406
rect 12728 11558 12756 12786
rect 13004 12186 13032 12922
rect 13096 12850 13124 13330
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 13188 12730 13216 14962
rect 13266 14240 13322 14249
rect 13266 14175 13322 14184
rect 12820 12158 13032 12186
rect 13096 12702 13216 12730
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12820 11150 12848 12158
rect 12992 12096 13044 12102
rect 12990 12064 12992 12073
rect 13044 12064 13046 12073
rect 12990 11999 13046 12008
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12912 11393 12940 11698
rect 13096 11676 13124 12702
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 13188 12238 13216 12582
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13280 12170 13308 14175
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13372 13190 13400 13874
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13372 12753 13400 12786
rect 13358 12744 13414 12753
rect 13358 12679 13414 12688
rect 13464 12628 13492 13874
rect 13648 12730 13676 15982
rect 13740 14958 13768 16050
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13740 14482 13768 14894
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 14292 14414 14320 16186
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13740 12850 13768 13126
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13648 12702 13768 12730
rect 13372 12600 13492 12628
rect 13372 12481 13400 12600
rect 13358 12472 13414 12481
rect 13358 12407 13414 12416
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 13176 11688 13228 11694
rect 13096 11648 13176 11676
rect 13176 11630 13228 11636
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 12898 11384 12954 11393
rect 12898 11319 12954 11328
rect 12992 11348 13044 11354
rect 12808 11144 12860 11150
rect 12806 11112 12808 11121
rect 12860 11112 12862 11121
rect 12806 11047 12862 11056
rect 12624 11008 12676 11014
rect 12530 10976 12586 10985
rect 12624 10950 12676 10956
rect 12530 10911 12586 10920
rect 12438 10160 12494 10169
rect 12438 10095 12494 10104
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12452 9654 12480 9862
rect 12544 9654 12572 10911
rect 12636 10826 12664 10950
rect 12636 10810 12848 10826
rect 12636 10804 12860 10810
rect 12636 10798 12808 10804
rect 12808 10746 12860 10752
rect 12624 10736 12676 10742
rect 12912 10690 12940 11319
rect 12992 11290 13044 11296
rect 13004 10713 13032 11290
rect 13096 10742 13124 11494
rect 13084 10736 13136 10742
rect 12624 10678 12676 10684
rect 12636 10062 12664 10678
rect 12820 10662 12940 10690
rect 12990 10704 13046 10713
rect 12714 10568 12770 10577
rect 12714 10503 12770 10512
rect 12728 10470 12756 10503
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12532 9512 12584 9518
rect 12636 9500 12664 9658
rect 12714 9616 12770 9625
rect 12714 9551 12770 9560
rect 12728 9518 12756 9551
rect 12584 9472 12664 9500
rect 12716 9512 12768 9518
rect 12532 9454 12584 9460
rect 12716 9454 12768 9460
rect 12716 9376 12768 9382
rect 12438 9344 12494 9353
rect 12716 9318 12768 9324
rect 12438 9279 12494 9288
rect 12452 8498 12480 9279
rect 12728 9110 12756 9318
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12440 8016 12492 8022
rect 12440 7958 12492 7964
rect 12452 7410 12480 7958
rect 12544 7585 12572 8774
rect 12820 8566 12848 10662
rect 13084 10678 13136 10684
rect 12990 10639 13046 10648
rect 12900 10464 12952 10470
rect 13096 10441 13124 10678
rect 12900 10406 12952 10412
rect 13082 10432 13138 10441
rect 12912 9466 12940 10406
rect 13082 10367 13138 10376
rect 13188 10305 13216 11630
rect 13280 10713 13308 12106
rect 13266 10704 13322 10713
rect 13266 10639 13322 10648
rect 13174 10296 13230 10305
rect 13174 10231 13230 10240
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 13004 9568 13032 10066
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 13096 9722 13124 9998
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13004 9540 13124 9568
rect 12912 9438 13032 9466
rect 13096 9450 13124 9540
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12636 7886 12664 8230
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12530 7576 12586 7585
rect 12530 7511 12586 7520
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 11992 5710 12020 6054
rect 12162 5944 12218 5953
rect 12162 5879 12218 5888
rect 12072 5840 12124 5846
rect 12070 5808 12072 5817
rect 12124 5808 12126 5817
rect 12070 5743 12126 5752
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11992 5001 12020 5646
rect 11978 4992 12034 5001
rect 11978 4927 12034 4936
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11992 4282 12020 4422
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 12084 4146 12112 5743
rect 12176 4146 12204 5879
rect 12268 5234 12296 6054
rect 12360 5914 12388 6190
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12452 5710 12480 7346
rect 12544 6322 12572 7511
rect 12622 7440 12678 7449
rect 12622 7375 12624 7384
rect 12676 7375 12678 7384
rect 12624 7346 12676 7352
rect 12728 7002 12756 7686
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12820 7177 12848 7278
rect 12806 7168 12862 7177
rect 12806 7103 12862 7112
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12440 5704 12492 5710
rect 12492 5664 12664 5692
rect 12440 5646 12492 5652
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12440 5024 12492 5030
rect 12544 5012 12572 5170
rect 12492 4984 12572 5012
rect 12440 4966 12492 4972
rect 12360 4826 12388 4966
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12636 4078 12664 5664
rect 12728 5234 12756 6938
rect 12912 5574 12940 9318
rect 13004 7410 13032 9438
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 13096 8838 13124 9386
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 13188 8022 13216 10134
rect 13372 9722 13400 12174
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13372 9353 13400 9522
rect 13358 9344 13414 9353
rect 13358 9279 13414 9288
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13280 8430 13308 8570
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13176 8016 13228 8022
rect 13176 7958 13228 7964
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 13188 7410 13216 7686
rect 12992 7404 13044 7410
rect 13176 7404 13228 7410
rect 13044 7364 13124 7392
rect 12992 7346 13044 7352
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 13004 5681 13032 6054
rect 13096 5846 13124 7364
rect 13176 7346 13228 7352
rect 13372 7274 13400 8298
rect 13360 7268 13412 7274
rect 13360 7210 13412 7216
rect 13266 7168 13322 7177
rect 13266 7103 13322 7112
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13188 5914 13216 6258
rect 13280 5914 13308 7103
rect 13372 6497 13400 7210
rect 13358 6488 13414 6497
rect 13358 6423 13414 6432
rect 13464 6322 13492 12378
rect 13740 12374 13768 12702
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13556 11898 13584 12174
rect 13832 11914 13860 13262
rect 13924 12730 13952 14350
rect 14292 13954 14320 14350
rect 14372 14340 14424 14346
rect 14372 14282 14424 14288
rect 14464 14340 14516 14346
rect 14464 14282 14516 14288
rect 14384 14074 14412 14282
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14292 13938 14412 13954
rect 14292 13932 14424 13938
rect 14292 13926 14372 13932
rect 14372 13874 14424 13880
rect 14188 13864 14240 13870
rect 14108 13824 14188 13852
rect 13924 12702 14044 12730
rect 14016 12646 14044 12702
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 14004 12640 14056 12646
rect 14108 12617 14136 13824
rect 14476 13818 14504 14282
rect 14240 13812 14504 13818
rect 14188 13806 14504 13812
rect 14200 13790 14504 13806
rect 14568 13818 14596 14894
rect 14660 13938 14688 17002
rect 14832 16516 14884 16522
rect 14832 16458 14884 16464
rect 14844 14414 14872 16458
rect 14936 15502 14964 17478
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15120 16794 15148 17138
rect 15108 16788 15160 16794
rect 15108 16730 15160 16736
rect 15016 16720 15068 16726
rect 15016 16662 15068 16668
rect 14924 15496 14976 15502
rect 14922 15464 14924 15473
rect 14976 15464 14978 15473
rect 15028 15434 15056 16662
rect 14922 15399 14978 15408
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 15120 14521 15148 16730
rect 15212 15162 15240 17138
rect 16040 17066 16068 17546
rect 16028 17060 16080 17066
rect 16028 17002 16080 17008
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15856 16250 15884 16594
rect 16040 16590 16068 17002
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16224 16590 16252 16934
rect 16500 16590 16528 18294
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16592 17678 16620 18226
rect 16684 17882 16712 18634
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16592 16590 16620 17614
rect 16776 17270 16804 18090
rect 16764 17264 16816 17270
rect 16764 17206 16816 17212
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 16488 16176 16540 16182
rect 16488 16118 16540 16124
rect 16500 16017 16528 16118
rect 16592 16114 16620 16526
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16486 16008 16542 16017
rect 16486 15943 16542 15952
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15106 14512 15162 14521
rect 15106 14447 15162 14456
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 15016 14408 15068 14414
rect 15068 14356 15148 14362
rect 15016 14350 15148 14356
rect 14844 14006 14872 14350
rect 15028 14334 15148 14350
rect 14832 14000 14884 14006
rect 14832 13942 14884 13948
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14844 13870 14872 13942
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14832 13864 14884 13870
rect 14568 13790 14688 13818
rect 14832 13806 14884 13812
rect 14554 13424 14610 13433
rect 14554 13359 14610 13368
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14292 12850 14320 13194
rect 14568 12918 14596 13359
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14004 12582 14056 12588
rect 14094 12608 14150 12617
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13648 11886 13860 11914
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13556 7886 13584 11018
rect 13648 11014 13676 11886
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13740 11529 13768 11766
rect 13820 11552 13872 11558
rect 13726 11520 13782 11529
rect 13820 11494 13872 11500
rect 13726 11455 13782 11464
rect 13832 11150 13860 11494
rect 13924 11150 13952 12582
rect 14094 12543 14150 12552
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14108 11150 14136 11698
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13648 10470 13676 10950
rect 13832 10742 13860 11086
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 14002 10704 14058 10713
rect 14002 10639 14004 10648
rect 14056 10639 14058 10648
rect 14004 10610 14056 10616
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13648 9110 13676 9998
rect 14016 9602 14044 10066
rect 13832 9592 14044 9602
rect 13832 9586 14056 9592
rect 13832 9574 14004 9586
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13648 8498 13676 8570
rect 13740 8498 13768 9318
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13740 8090 13768 8230
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13636 7948 13688 7954
rect 13688 7908 13768 7936
rect 13636 7890 13688 7896
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13556 6662 13584 7346
rect 13648 7002 13676 7346
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13740 6322 13768 7908
rect 13832 6798 13860 9574
rect 14004 9528 14056 9534
rect 14004 9104 14056 9110
rect 14004 9046 14056 9052
rect 14016 8430 14044 9046
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13924 7410 13952 8230
rect 14016 7993 14044 8366
rect 14002 7984 14058 7993
rect 14002 7919 14058 7928
rect 14016 7410 14044 7919
rect 14108 7886 14136 10406
rect 14200 8922 14228 12310
rect 14292 11506 14320 12786
rect 14476 12753 14504 12786
rect 14462 12744 14518 12753
rect 14462 12679 14518 12688
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14476 12238 14504 12582
rect 14568 12374 14596 12854
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14372 12232 14424 12238
rect 14370 12200 14372 12209
rect 14464 12232 14516 12238
rect 14424 12200 14426 12209
rect 14464 12174 14516 12180
rect 14370 12135 14426 12144
rect 14384 11626 14412 12135
rect 14660 12102 14688 13790
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14752 12850 14780 13262
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14844 12714 14872 13670
rect 14832 12708 14884 12714
rect 14832 12650 14884 12656
rect 14830 12608 14886 12617
rect 14830 12543 14886 12552
rect 14844 12434 14872 12543
rect 14752 12406 14872 12434
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14476 11762 14504 12038
rect 14660 11898 14688 12038
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14372 11620 14424 11626
rect 14372 11562 14424 11568
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14292 11478 14412 11506
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 10674 14320 10950
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14384 10452 14412 11478
rect 14568 11354 14596 11562
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 14476 10577 14504 11222
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14462 10568 14518 10577
rect 14462 10503 14518 10512
rect 14568 10452 14596 11154
rect 14660 11132 14688 11698
rect 14752 11286 14780 12406
rect 14830 12336 14886 12345
rect 14830 12271 14886 12280
rect 14844 12238 14872 12271
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14740 11280 14792 11286
rect 14740 11222 14792 11228
rect 14660 11104 14780 11132
rect 14752 10470 14780 11104
rect 14384 10424 14596 10452
rect 14568 10266 14596 10424
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 14278 9616 14334 9625
rect 14384 9586 14412 9930
rect 14568 9722 14596 10066
rect 14752 10062 14780 10406
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14278 9551 14280 9560
rect 14332 9551 14334 9560
rect 14372 9580 14424 9586
rect 14280 9522 14332 9528
rect 14372 9522 14424 9528
rect 14476 9450 14504 9658
rect 14752 9586 14780 9998
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14476 9058 14504 9114
rect 14292 9042 14504 9058
rect 14280 9036 14504 9042
rect 14332 9030 14504 9036
rect 14280 8978 14332 8984
rect 14464 8968 14516 8974
rect 14200 8894 14320 8922
rect 14464 8910 14516 8916
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14200 8090 14228 8774
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13084 5840 13136 5846
rect 13084 5782 13136 5788
rect 13634 5808 13690 5817
rect 13544 5772 13596 5778
rect 13634 5743 13690 5752
rect 13544 5714 13596 5720
rect 12990 5672 13046 5681
rect 12990 5607 13046 5616
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 13556 5234 13584 5714
rect 13648 5710 13676 5743
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 12992 5024 13044 5030
rect 12912 4984 12992 5012
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 12084 3194 12112 3470
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12544 3194 12572 3334
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12912 3126 12940 4984
rect 12992 4966 13044 4972
rect 13096 4282 13124 5170
rect 13648 5166 13676 5510
rect 13740 5166 13768 6258
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13832 5370 13860 5510
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13912 5024 13964 5030
rect 13634 4992 13690 5001
rect 13912 4966 13964 4972
rect 13634 4927 13690 4936
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13280 4622 13308 4694
rect 13464 4622 13492 4762
rect 13648 4690 13676 4927
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13268 4616 13320 4622
rect 13174 4584 13230 4593
rect 13268 4558 13320 4564
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13174 4519 13230 4528
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 13188 4128 13216 4519
rect 13280 4282 13308 4558
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13372 4214 13400 4422
rect 13360 4208 13412 4214
rect 13360 4150 13412 4156
rect 13268 4140 13320 4146
rect 13188 4100 13268 4128
rect 13268 4082 13320 4088
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13266 4040 13322 4049
rect 13266 3975 13322 3984
rect 13082 3632 13138 3641
rect 13082 3567 13138 3576
rect 13096 3534 13124 3567
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12716 3120 12768 3126
rect 12714 3088 12716 3097
rect 12900 3120 12952 3126
rect 12768 3088 12770 3097
rect 12900 3062 12952 3068
rect 12714 3023 12770 3032
rect 13280 2990 13308 3975
rect 13556 3670 13584 4082
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13464 3194 13492 3470
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13556 3058 13584 3606
rect 13648 3466 13676 4626
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13740 3913 13768 4082
rect 13726 3904 13782 3913
rect 13726 3839 13782 3848
rect 13832 3738 13860 4558
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13924 2922 13952 4966
rect 14108 4554 14136 7482
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14200 5302 14228 7346
rect 14292 7002 14320 8894
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14384 8566 14412 8774
rect 14476 8634 14504 8910
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 14372 8424 14424 8430
rect 14370 8392 14372 8401
rect 14424 8392 14426 8401
rect 14370 8327 14426 8336
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14384 6390 14412 7142
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14568 6746 14596 9522
rect 14660 8537 14688 9522
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14752 8634 14780 8910
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14646 8528 14702 8537
rect 14844 8498 14872 12038
rect 14936 10810 14964 13874
rect 15120 13802 15148 14334
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 15016 13456 15068 13462
rect 15016 13398 15068 13404
rect 15028 13326 15056 13398
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 15028 12918 15056 13126
rect 15016 12912 15068 12918
rect 15016 12854 15068 12860
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 15028 12209 15056 12650
rect 15014 12200 15070 12209
rect 15014 12135 15070 12144
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 15028 11558 15056 12038
rect 15016 11552 15068 11558
rect 15014 11520 15016 11529
rect 15068 11520 15070 11529
rect 15014 11455 15070 11464
rect 15028 11150 15056 11455
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 14922 10704 14978 10713
rect 14922 10639 14978 10648
rect 14936 9586 14964 10639
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 15028 9518 15056 10950
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 14924 8968 14976 8974
rect 14922 8936 14924 8945
rect 14976 8936 14978 8945
rect 14922 8871 14978 8880
rect 14922 8800 14978 8809
rect 14922 8735 14978 8744
rect 14646 8463 14702 8472
rect 14832 8492 14884 8498
rect 14660 8362 14688 8463
rect 14832 8434 14884 8440
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14660 7478 14688 7754
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 14752 7342 14780 8230
rect 14740 7336 14792 7342
rect 14740 7278 14792 7284
rect 14830 7304 14886 7313
rect 14830 7239 14886 7248
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14372 6384 14424 6390
rect 14278 6352 14334 6361
rect 14372 6326 14424 6332
rect 14278 6287 14280 6296
rect 14332 6287 14334 6296
rect 14280 6258 14332 6264
rect 14476 6118 14504 6734
rect 14568 6718 14688 6746
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 6322 14596 6598
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14556 6180 14608 6186
rect 14556 6122 14608 6128
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14370 5672 14426 5681
rect 14370 5607 14372 5616
rect 14424 5607 14426 5616
rect 14372 5578 14424 5584
rect 14278 5536 14334 5545
rect 14278 5471 14334 5480
rect 14188 5296 14240 5302
rect 14188 5238 14240 5244
rect 14292 5234 14320 5471
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14476 4758 14504 6054
rect 14568 5370 14596 6122
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14464 4752 14516 4758
rect 14464 4694 14516 4700
rect 14096 4548 14148 4554
rect 14096 4490 14148 4496
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14200 4078 14228 4422
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 14292 3670 14320 4014
rect 14280 3664 14332 3670
rect 14280 3606 14332 3612
rect 14384 3534 14412 4082
rect 14568 3534 14596 5306
rect 14660 4010 14688 6718
rect 14752 4758 14780 7142
rect 14844 4826 14872 7239
rect 14936 6798 14964 8735
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 14936 6186 14964 6734
rect 14924 6180 14976 6186
rect 14924 6122 14976 6128
rect 14922 5944 14978 5953
rect 14922 5879 14978 5888
rect 14936 5710 14964 5879
rect 14924 5704 14976 5710
rect 15028 5692 15056 9454
rect 15120 7546 15148 13738
rect 15212 13240 15240 15098
rect 15488 14822 15516 15098
rect 15764 15026 15792 15642
rect 16118 15600 16174 15609
rect 16118 15535 16174 15544
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15488 14414 15516 14758
rect 15672 14482 15700 14758
rect 15764 14482 15792 14962
rect 15948 14634 15976 15302
rect 15948 14606 16068 14634
rect 15936 14544 15988 14550
rect 15936 14486 15988 14492
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15304 13530 15332 14350
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15488 14006 15516 14214
rect 15476 14000 15528 14006
rect 15476 13942 15528 13948
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15292 13252 15344 13258
rect 15212 13212 15292 13240
rect 15292 13194 15344 13200
rect 15396 13138 15424 13874
rect 15212 13110 15424 13138
rect 15212 12442 15240 13110
rect 15580 13002 15608 14418
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15672 13326 15700 13806
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 15396 12974 15608 13002
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15198 11792 15254 11801
rect 15198 11727 15254 11736
rect 15212 11354 15240 11727
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15212 10606 15240 10950
rect 15304 10674 15332 12038
rect 15396 11098 15424 12974
rect 15672 12374 15700 13126
rect 15764 12850 15792 13330
rect 15948 13326 15976 14486
rect 16040 13870 16068 14606
rect 16028 13864 16080 13870
rect 16026 13832 16028 13841
rect 16080 13832 16082 13841
rect 16026 13767 16082 13776
rect 16132 13530 16160 15535
rect 16304 14884 16356 14890
rect 16304 14826 16356 14832
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15660 12368 15712 12374
rect 15474 12336 15530 12345
rect 15660 12310 15712 12316
rect 15474 12271 15530 12280
rect 15488 11218 15516 12271
rect 15566 11928 15622 11937
rect 15566 11863 15622 11872
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15396 11070 15516 11098
rect 15580 11082 15608 11863
rect 15672 11558 15700 12310
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15764 11336 15792 12786
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15856 11626 15884 12582
rect 15948 12442 15976 13262
rect 16132 12850 16160 13466
rect 16316 12850 16344 14826
rect 16500 14550 16528 15943
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16684 15502 16712 15846
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16580 15360 16632 15366
rect 16776 15314 16804 16390
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 16580 15302 16632 15308
rect 16488 14544 16540 14550
rect 16488 14486 16540 14492
rect 16592 13938 16620 15302
rect 16684 15286 16804 15314
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16408 12918 16436 13126
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16120 12844 16172 12850
rect 16040 12804 16120 12832
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15764 11308 15884 11336
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15488 11014 15516 11070
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15580 10810 15608 11018
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15566 10704 15622 10713
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15476 10668 15528 10674
rect 15566 10639 15568 10648
rect 15476 10610 15528 10616
rect 15620 10639 15622 10648
rect 15568 10610 15620 10616
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15488 10062 15516 10610
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 15212 9450 15240 9930
rect 15200 9444 15252 9450
rect 15200 9386 15252 9392
rect 15212 8498 15240 9386
rect 15396 9382 15424 9998
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15292 9104 15344 9110
rect 15292 9046 15344 9052
rect 15304 8498 15332 9046
rect 15488 8786 15516 9998
rect 15396 8758 15516 8786
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15304 8022 15332 8434
rect 15292 8016 15344 8022
rect 15292 7958 15344 7964
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15304 7410 15332 7686
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15200 7336 15252 7342
rect 15198 7304 15200 7313
rect 15252 7304 15254 7313
rect 15198 7239 15254 7248
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15108 6792 15160 6798
rect 15212 6780 15240 7142
rect 15290 6896 15346 6905
rect 15290 6831 15346 6840
rect 15304 6798 15332 6831
rect 15160 6752 15240 6780
rect 15108 6734 15160 6740
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15120 5710 15148 5850
rect 14976 5664 15056 5692
rect 14924 5646 14976 5652
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14740 4752 14792 4758
rect 14740 4694 14792 4700
rect 15028 4214 15056 5664
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15212 5642 15240 6752
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15200 5636 15252 5642
rect 15200 5578 15252 5584
rect 15212 5098 15240 5578
rect 15304 5234 15332 6190
rect 15396 5710 15424 8758
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15488 7886 15516 8570
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15488 6798 15516 7822
rect 15580 7206 15608 10610
rect 15672 8974 15700 11086
rect 15764 10674 15792 11154
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15764 10266 15792 10610
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15856 10062 15884 11308
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15948 9908 15976 11494
rect 16040 10674 16068 12804
rect 16120 12786 16172 12792
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16224 12306 16252 12582
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16224 11082 16252 12242
rect 16212 11076 16264 11082
rect 16212 11018 16264 11024
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 16132 10538 16160 10950
rect 16120 10532 16172 10538
rect 16120 10474 16172 10480
rect 16316 10266 16344 12786
rect 16396 12708 16448 12714
rect 16396 12650 16448 12656
rect 16408 12170 16436 12650
rect 16396 12164 16448 12170
rect 16396 12106 16448 12112
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16304 10260 16356 10266
rect 16304 10202 16356 10208
rect 16028 9920 16080 9926
rect 15948 9880 16028 9908
rect 16028 9862 16080 9868
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15660 8832 15712 8838
rect 15658 8800 15660 8809
rect 15712 8800 15714 8809
rect 15658 8735 15714 8744
rect 15750 8528 15806 8537
rect 15856 8498 15884 9454
rect 15948 9110 15976 9454
rect 15936 9104 15988 9110
rect 15936 9046 15988 9052
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15948 8566 15976 8774
rect 15936 8560 15988 8566
rect 15936 8502 15988 8508
rect 15750 8463 15752 8472
rect 15804 8463 15806 8472
rect 15844 8492 15896 8498
rect 15752 8434 15804 8440
rect 15844 8434 15896 8440
rect 15764 8294 15792 8434
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15672 6458 15700 8026
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15764 7410 15792 7958
rect 15856 7750 15884 8434
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15764 6322 15792 6938
rect 15856 6934 15884 7686
rect 15844 6928 15896 6934
rect 15844 6870 15896 6876
rect 15856 6458 15884 6870
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15936 6384 15988 6390
rect 15936 6326 15988 6332
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15764 5914 15792 6258
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15488 5302 15516 5510
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15476 5296 15528 5302
rect 15476 5238 15528 5244
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15200 5092 15252 5098
rect 15200 5034 15252 5040
rect 15016 4208 15068 4214
rect 15016 4150 15068 4156
rect 15212 4146 15240 5034
rect 15764 4826 15792 5306
rect 15948 4826 15976 6326
rect 16040 5302 16068 9862
rect 16120 9648 16172 9654
rect 16120 9590 16172 9596
rect 16132 9353 16160 9590
rect 16118 9344 16174 9353
rect 16118 9279 16174 9288
rect 16118 9072 16174 9081
rect 16118 9007 16174 9016
rect 16132 8974 16160 9007
rect 16224 8974 16252 10202
rect 16408 9994 16436 10610
rect 16578 10432 16634 10441
rect 16578 10367 16634 10376
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 16486 9616 16542 9625
rect 16486 9551 16542 9560
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16408 8974 16436 9318
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16132 8634 16160 8910
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16132 8090 16160 8434
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16224 7886 16252 8910
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16224 6866 16252 7346
rect 16408 7342 16436 8910
rect 16500 8498 16528 9551
rect 16592 8650 16620 10367
rect 16684 9586 16712 15286
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16776 13870 16804 14010
rect 16868 13954 16896 15438
rect 17052 15162 17080 16050
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 17144 15026 17172 15846
rect 17776 15632 17828 15638
rect 17222 15600 17278 15609
rect 17776 15574 17828 15580
rect 17222 15535 17224 15544
rect 17276 15535 17278 15544
rect 17224 15506 17276 15512
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 16960 14074 16988 14962
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 17052 14074 17080 14214
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 17040 14068 17092 14074
rect 17040 14010 17092 14016
rect 16868 13926 16988 13954
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16776 11665 16804 11698
rect 16762 11656 16818 11665
rect 16960 11626 16988 13926
rect 16762 11591 16818 11600
rect 16948 11620 17000 11626
rect 16948 11562 17000 11568
rect 17144 10742 17172 14962
rect 17236 12850 17264 15098
rect 17512 14890 17540 15438
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 17500 14340 17552 14346
rect 17500 14282 17552 14288
rect 17328 12986 17356 14282
rect 17512 14074 17540 14282
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17604 13938 17632 15302
rect 17788 14482 17816 15574
rect 18052 15088 18104 15094
rect 17958 15056 18014 15065
rect 18052 15030 18104 15036
rect 17958 14991 17960 15000
rect 18012 14991 18014 15000
rect 17960 14962 18012 14968
rect 17684 14476 17736 14482
rect 17684 14418 17736 14424
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17696 13938 17724 14418
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17420 13462 17448 13874
rect 17604 13841 17632 13874
rect 17590 13832 17646 13841
rect 17590 13767 17646 13776
rect 17788 13530 17816 14418
rect 17958 14376 18014 14385
rect 17958 14311 18014 14320
rect 17972 14074 18000 14311
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18064 13705 18092 15030
rect 18050 13696 18106 13705
rect 18050 13631 18106 13640
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17408 13456 17460 13462
rect 17408 13398 17460 13404
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 17222 11248 17278 11257
rect 17222 11183 17278 11192
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 17052 10198 17080 10542
rect 17144 10470 17172 10678
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17040 10192 17092 10198
rect 17040 10134 17092 10140
rect 17236 10062 17264 11183
rect 17328 10810 17356 12106
rect 17512 11082 17540 12582
rect 17788 12434 17816 13466
rect 17696 12406 17816 12434
rect 17696 12238 17724 12406
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17592 11620 17644 11626
rect 17592 11562 17644 11568
rect 17500 11076 17552 11082
rect 17500 11018 17552 11024
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17408 10736 17460 10742
rect 17408 10678 17460 10684
rect 17224 10056 17276 10062
rect 17224 9998 17276 10004
rect 16948 9988 17000 9994
rect 16948 9930 17000 9936
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16592 8622 16712 8650
rect 16580 8560 16632 8566
rect 16580 8502 16632 8508
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15672 4146 15700 4626
rect 16132 4554 16160 5714
rect 16224 5234 16252 6394
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16120 4548 16172 4554
rect 16120 4490 16172 4496
rect 16132 4214 16160 4490
rect 16224 4282 16252 5170
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16316 4622 16344 5102
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16120 4208 16172 4214
rect 16120 4150 16172 4156
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 14648 4004 14700 4010
rect 14648 3946 14700 3952
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14660 3466 14688 3946
rect 15672 3602 15700 4082
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 16132 3534 16160 4150
rect 16316 4146 16344 4558
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16592 3942 16620 8502
rect 16684 5574 16712 8622
rect 16868 7342 16896 9114
rect 16960 8498 16988 9930
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 17052 8974 17080 9318
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 17052 8566 17080 8910
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16960 7410 16988 8434
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16868 6934 16896 7278
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 16868 6322 16896 6870
rect 16948 6724 17000 6730
rect 16948 6666 17000 6672
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16868 5778 16896 6258
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16684 5370 16712 5510
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16776 4010 16804 5578
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 16960 3942 16988 6666
rect 17052 6390 17080 8502
rect 17236 6458 17264 9998
rect 17420 8974 17448 10678
rect 17604 10538 17632 11562
rect 17696 11218 17724 12174
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17972 11354 18000 11698
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17592 10532 17644 10538
rect 17592 10474 17644 10480
rect 17604 9674 17632 10474
rect 17604 9646 17724 9674
rect 17696 9586 17724 9646
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 17052 6254 17080 6326
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 17420 5710 17448 8910
rect 17696 6730 17724 9522
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17972 7585 18000 7686
rect 17958 7576 18014 7585
rect 17958 7511 18014 7520
rect 17684 6724 17736 6730
rect 17684 6666 17736 6672
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 14648 3460 14700 3466
rect 14648 3402 14700 3408
rect 15396 3194 15424 3470
rect 16592 3466 16620 3878
rect 16580 3460 16632 3466
rect 16580 3402 16632 3408
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 13004 2446 13032 2790
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 6472 800 6500 2246
rect 9048 800 9076 2246
rect 9692 800 9720 2246
rect 13556 800 13584 2246
rect 6458 0 6514 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 13542 0 13598 800
<< via2 >>
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 3054 16108 3110 16144
rect 3054 16088 3056 16108
rect 3056 16088 3108 16108
rect 3108 16088 3110 16108
rect 2962 15544 3018 15600
rect 846 14492 848 14512
rect 848 14492 900 14512
rect 900 14492 902 14512
rect 846 14456 902 14492
rect 1490 13676 1492 13696
rect 1492 13676 1544 13696
rect 1544 13676 1546 13696
rect 1490 13640 1546 13676
rect 1030 8880 1086 8936
rect 1490 5516 1492 5536
rect 1492 5516 1544 5536
rect 1544 5516 1546 5536
rect 1490 5480 1546 5516
rect 2502 13368 2558 13424
rect 3238 14900 3240 14920
rect 3240 14900 3292 14920
rect 3292 14900 3294 14920
rect 2870 13268 2872 13288
rect 2872 13268 2924 13288
rect 2924 13268 2926 13288
rect 2870 13232 2926 13268
rect 2778 13096 2834 13152
rect 3238 14864 3294 14900
rect 3146 13268 3148 13288
rect 3148 13268 3200 13288
rect 3200 13268 3202 13288
rect 3146 13232 3202 13268
rect 3054 12552 3110 12608
rect 2594 11092 2596 11112
rect 2596 11092 2648 11112
rect 2648 11092 2650 11112
rect 2594 11056 2650 11092
rect 3514 15000 3570 15056
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4618 15408 4674 15464
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 5354 16496 5410 16552
rect 5262 16088 5318 16144
rect 5078 15988 5080 16008
rect 5080 15988 5132 16008
rect 5132 15988 5134 16008
rect 5078 15952 5134 15988
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4066 13812 4068 13832
rect 4068 13812 4120 13832
rect 4120 13812 4122 13832
rect 4066 13776 4122 13812
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 5078 15428 5134 15464
rect 5078 15408 5080 15428
rect 5080 15408 5132 15428
rect 5132 15408 5134 15428
rect 5538 15952 5594 16008
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4710 14356 4712 14376
rect 4712 14356 4764 14376
rect 4764 14356 4766 14376
rect 4710 14320 4766 14356
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4526 12144 4582 12200
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4894 13524 4950 13560
rect 4894 13504 4896 13524
rect 4896 13504 4948 13524
rect 4948 13504 4950 13524
rect 5538 15000 5594 15056
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4894 12688 4950 12744
rect 5078 12416 5134 12472
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 5078 11736 5134 11792
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 3054 9580 3110 9616
rect 3054 9560 3056 9580
rect 3056 9560 3108 9580
rect 3108 9560 3110 9580
rect 2962 9016 3018 9072
rect 2778 8744 2834 8800
rect 3146 8472 3202 8528
rect 3330 9696 3386 9752
rect 4066 10512 4122 10568
rect 3882 10104 3938 10160
rect 3054 5616 3110 5672
rect 3790 8744 3846 8800
rect 3790 8472 3846 8528
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4434 10104 4490 10160
rect 6366 16088 6422 16144
rect 6090 15428 6146 15464
rect 6090 15408 6092 15428
rect 6092 15408 6144 15428
rect 6144 15408 6146 15428
rect 5722 13948 5724 13968
rect 5724 13948 5776 13968
rect 5776 13948 5778 13968
rect 5722 13912 5778 13948
rect 5722 13232 5778 13288
rect 4986 10512 5042 10568
rect 4710 9968 4766 10024
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4434 9016 4490 9072
rect 4158 8916 4160 8936
rect 4160 8916 4212 8936
rect 4212 8916 4214 8936
rect 4158 8880 4214 8916
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 3514 6316 3570 6352
rect 3514 6296 3516 6316
rect 3516 6296 3568 6316
rect 3568 6296 3570 6316
rect 3698 6296 3754 6352
rect 3606 5752 3662 5808
rect 2778 3440 2834 3496
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 5262 9968 5318 10024
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 5262 9632 5318 9688
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 5170 8492 5226 8528
rect 5170 8472 5172 8492
rect 5172 8472 5224 8492
rect 5224 8472 5226 8492
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 5998 12824 6054 12880
rect 6274 15408 6330 15464
rect 6182 14184 6238 14240
rect 6182 13776 6238 13832
rect 6458 15408 6514 15464
rect 6826 14764 6828 14784
rect 6828 14764 6880 14784
rect 6880 14764 6882 14784
rect 6826 14728 6882 14764
rect 5906 10512 5962 10568
rect 5814 10376 5870 10432
rect 6090 11076 6146 11112
rect 6090 11056 6092 11076
rect 6092 11056 6144 11076
rect 6144 11056 6146 11076
rect 5354 7284 5356 7304
rect 5356 7284 5408 7304
rect 5408 7284 5410 7304
rect 5354 7248 5410 7284
rect 4894 6296 4950 6352
rect 4802 6160 4858 6216
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 5722 9832 5778 9888
rect 5906 9580 5962 9616
rect 5906 9560 5908 9580
rect 5908 9560 5960 9580
rect 5960 9560 5962 9580
rect 5814 9424 5870 9480
rect 5998 8508 6000 8528
rect 6000 8508 6052 8528
rect 6052 8508 6054 8528
rect 5998 8472 6054 8508
rect 6918 14184 6974 14240
rect 6918 13776 6974 13832
rect 7194 13524 7250 13560
rect 7194 13504 7196 13524
rect 7196 13504 7248 13524
rect 7248 13504 7250 13524
rect 6918 12724 6920 12744
rect 6920 12724 6972 12744
rect 6972 12724 6974 12744
rect 6918 12688 6974 12724
rect 6458 9580 6514 9616
rect 6458 9560 6460 9580
rect 6460 9560 6512 9580
rect 6512 9560 6514 9580
rect 6642 9560 6698 9616
rect 6918 11192 6974 11248
rect 6826 11092 6828 11112
rect 6828 11092 6880 11112
rect 6880 11092 6882 11112
rect 6826 11056 6882 11092
rect 7746 15544 7802 15600
rect 7838 15408 7894 15464
rect 7102 10376 7158 10432
rect 5722 6740 5724 6760
rect 5724 6740 5776 6760
rect 5776 6740 5778 6760
rect 5722 6704 5778 6740
rect 5998 7828 6000 7848
rect 6000 7828 6052 7848
rect 6052 7828 6054 7848
rect 5998 7792 6054 7828
rect 5998 6976 6054 7032
rect 5354 4548 5410 4584
rect 5354 4528 5356 4548
rect 5356 4528 5408 4548
rect 5408 4528 5410 4548
rect 5906 5344 5962 5400
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 6918 9016 6974 9072
rect 6642 8472 6698 8528
rect 6550 7928 6606 7984
rect 6366 6976 6422 7032
rect 6458 6296 6514 6352
rect 6918 8744 6974 8800
rect 7562 9696 7618 9752
rect 7746 12552 7802 12608
rect 8206 15272 8262 15328
rect 8206 14728 8262 14784
rect 7930 11464 7986 11520
rect 8298 11620 8354 11656
rect 8298 11600 8300 11620
rect 8300 11600 8352 11620
rect 8352 11600 8354 11620
rect 7194 8336 7250 8392
rect 6918 5480 6974 5536
rect 7286 8200 7342 8256
rect 7378 5888 7434 5944
rect 7010 3984 7066 4040
rect 6366 2896 6422 2952
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 7654 8336 7710 8392
rect 7654 7928 7710 7984
rect 8114 9016 8170 9072
rect 7930 6840 7986 6896
rect 7562 6432 7618 6488
rect 7838 6432 7894 6488
rect 7746 5888 7802 5944
rect 8298 10512 8354 10568
rect 9862 17756 9864 17776
rect 9864 17756 9916 17776
rect 9916 17756 9918 17776
rect 9862 17720 9918 17756
rect 10506 17720 10562 17776
rect 8758 16224 8814 16280
rect 8574 15544 8630 15600
rect 8574 14320 8630 14376
rect 8942 15852 8944 15872
rect 8944 15852 8996 15872
rect 8996 15852 8998 15872
rect 8942 15816 8998 15852
rect 8942 15544 8998 15600
rect 8574 13268 8576 13288
rect 8576 13268 8628 13288
rect 8628 13268 8630 13288
rect 8574 13232 8630 13268
rect 8574 12280 8630 12336
rect 8574 12008 8630 12064
rect 8758 10920 8814 10976
rect 8758 10668 8814 10704
rect 8758 10648 8760 10668
rect 8760 10648 8812 10668
rect 8812 10648 8814 10668
rect 8666 10412 8668 10432
rect 8668 10412 8720 10432
rect 8720 10412 8722 10432
rect 8666 10376 8722 10412
rect 9678 16632 9734 16688
rect 9310 15952 9366 16008
rect 9586 16088 9642 16144
rect 9310 15428 9366 15464
rect 9586 15816 9642 15872
rect 9862 16088 9918 16144
rect 9954 15816 10010 15872
rect 9310 15408 9312 15428
rect 9312 15408 9364 15428
rect 9364 15408 9366 15428
rect 9218 14864 9274 14920
rect 9586 15272 9642 15328
rect 9402 15036 9404 15056
rect 9404 15036 9456 15056
rect 9456 15036 9458 15056
rect 9402 15000 9458 15036
rect 9402 14864 9458 14920
rect 8942 12008 8998 12064
rect 9494 14320 9550 14376
rect 9678 14320 9734 14376
rect 9586 14048 9642 14104
rect 9126 11192 9182 11248
rect 9954 15408 10010 15464
rect 9954 14456 10010 14512
rect 9862 13932 9918 13968
rect 9862 13912 9864 13932
rect 9864 13912 9916 13932
rect 9916 13912 9918 13932
rect 9678 13504 9734 13560
rect 9770 13368 9826 13424
rect 9770 12960 9826 13016
rect 9494 12416 9550 12472
rect 9770 12416 9826 12472
rect 9218 10668 9274 10704
rect 9218 10648 9220 10668
rect 9220 10648 9272 10668
rect 9272 10648 9274 10668
rect 8574 10004 8576 10024
rect 8576 10004 8628 10024
rect 8628 10004 8630 10024
rect 8574 9968 8630 10004
rect 8574 9832 8630 9888
rect 8482 8608 8538 8664
rect 8298 8336 8354 8392
rect 8574 7792 8630 7848
rect 8482 5752 8538 5808
rect 8758 6160 8814 6216
rect 9034 8336 9090 8392
rect 9770 12008 9826 12064
rect 9862 11600 9918 11656
rect 9586 11464 9642 11520
rect 9770 11464 9826 11520
rect 9678 11328 9734 11384
rect 10046 11600 10102 11656
rect 9494 10260 9550 10296
rect 9494 10240 9496 10260
rect 9496 10240 9548 10260
rect 9548 10240 9550 10260
rect 9494 10004 9496 10024
rect 9496 10004 9548 10024
rect 9548 10004 9550 10024
rect 9494 9968 9550 10004
rect 9402 9832 9458 9888
rect 9218 7928 9274 7984
rect 8850 5344 8906 5400
rect 8850 5228 8906 5264
rect 8850 5208 8852 5228
rect 8852 5208 8904 5228
rect 8904 5208 8906 5228
rect 8666 3052 8722 3088
rect 8666 3032 8668 3052
rect 8668 3032 8720 3052
rect 8720 3032 8722 3052
rect 10230 15000 10286 15056
rect 10874 16632 10930 16688
rect 10414 13912 10470 13968
rect 10230 13776 10286 13832
rect 10414 13504 10470 13560
rect 10506 13368 10562 13424
rect 10690 12688 10746 12744
rect 10782 12416 10838 12472
rect 11334 15680 11390 15736
rect 11334 14184 11390 14240
rect 10230 11464 10286 11520
rect 10322 11328 10378 11384
rect 10138 10648 10194 10704
rect 9954 8336 10010 8392
rect 9586 6196 9588 6216
rect 9588 6196 9640 6216
rect 9640 6196 9642 6216
rect 9586 6160 9642 6196
rect 9494 5344 9550 5400
rect 10046 7384 10102 7440
rect 10230 8200 10286 8256
rect 10506 11328 10562 11384
rect 10598 9696 10654 9752
rect 10414 9288 10470 9344
rect 10322 7248 10378 7304
rect 11058 11872 11114 11928
rect 11334 13096 11390 13152
rect 11518 13096 11574 13152
rect 11242 12416 11298 12472
rect 11610 12552 11666 12608
rect 10874 10140 10876 10160
rect 10876 10140 10928 10160
rect 10928 10140 10930 10160
rect 10874 10104 10930 10140
rect 10414 6316 10470 6352
rect 10414 6296 10416 6316
rect 10416 6296 10468 6316
rect 10468 6296 10470 6316
rect 10322 5752 10378 5808
rect 9586 3848 9642 3904
rect 10690 7520 10746 7576
rect 11058 10648 11114 10704
rect 11334 10376 11390 10432
rect 11150 10240 11206 10296
rect 10874 8608 10930 8664
rect 10966 7112 11022 7168
rect 11518 10376 11574 10432
rect 11702 12280 11758 12336
rect 12070 16632 12126 16688
rect 12622 16224 12678 16280
rect 12898 16088 12954 16144
rect 12346 14456 12402 14512
rect 11886 12844 11942 12880
rect 11886 12824 11888 12844
rect 11888 12824 11940 12844
rect 11940 12824 11942 12844
rect 12346 12980 12402 13016
rect 12346 12960 12348 12980
rect 12348 12960 12400 12980
rect 12400 12960 12402 12980
rect 12254 11872 12310 11928
rect 11886 10784 11942 10840
rect 12070 11056 12126 11112
rect 12806 15036 12808 15056
rect 12808 15036 12860 15056
rect 12860 15036 12862 15056
rect 12806 15000 12862 15036
rect 13450 15544 13506 15600
rect 12990 13268 12992 13288
rect 12992 13268 13044 13288
rect 13044 13268 13046 13288
rect 12990 13232 13046 13268
rect 12530 12144 12586 12200
rect 12438 11600 12494 11656
rect 11794 10512 11850 10568
rect 11886 9696 11942 9752
rect 11518 9016 11574 9072
rect 11518 7964 11520 7984
rect 11520 7964 11572 7984
rect 11572 7964 11574 7984
rect 11518 7928 11574 7964
rect 10782 6432 10838 6488
rect 10598 5480 10654 5536
rect 11518 7248 11574 7304
rect 11334 6296 11390 6352
rect 10598 4120 10654 4176
rect 9954 3476 9956 3496
rect 9956 3476 10008 3496
rect 10008 3476 10010 3496
rect 9954 3440 10010 3476
rect 10690 3440 10746 3496
rect 11886 8608 11942 8664
rect 12254 9288 12310 9344
rect 12254 9016 12310 9072
rect 11794 6704 11850 6760
rect 12070 6840 12126 6896
rect 10322 2896 10378 2952
rect 13266 14184 13322 14240
rect 12990 12044 12992 12064
rect 12992 12044 13044 12064
rect 13044 12044 13046 12064
rect 12990 12008 13046 12044
rect 13358 12688 13414 12744
rect 13358 12416 13414 12472
rect 12898 11328 12954 11384
rect 12806 11092 12808 11112
rect 12808 11092 12860 11112
rect 12860 11092 12862 11112
rect 12806 11056 12862 11092
rect 12530 10920 12586 10976
rect 12438 10104 12494 10160
rect 12714 10512 12770 10568
rect 12714 9560 12770 9616
rect 12438 9288 12494 9344
rect 12990 10648 13046 10704
rect 13082 10376 13138 10432
rect 13266 10648 13322 10704
rect 13174 10240 13230 10296
rect 12530 7520 12586 7576
rect 12162 5888 12218 5944
rect 12070 5788 12072 5808
rect 12072 5788 12124 5808
rect 12124 5788 12126 5808
rect 12070 5752 12126 5788
rect 11978 4936 12034 4992
rect 12622 7404 12678 7440
rect 12622 7384 12624 7404
rect 12624 7384 12676 7404
rect 12676 7384 12678 7404
rect 12806 7112 12862 7168
rect 13358 9288 13414 9344
rect 13266 7112 13322 7168
rect 13358 6432 13414 6488
rect 14922 15444 14924 15464
rect 14924 15444 14976 15464
rect 14976 15444 14978 15464
rect 14922 15408 14978 15444
rect 16486 15952 16542 16008
rect 15106 14456 15162 14512
rect 14554 13368 14610 13424
rect 13726 11464 13782 11520
rect 14094 12552 14150 12608
rect 14002 10668 14058 10704
rect 14002 10648 14004 10668
rect 14004 10648 14056 10668
rect 14056 10648 14058 10668
rect 14002 7928 14058 7984
rect 14462 12688 14518 12744
rect 14370 12180 14372 12200
rect 14372 12180 14424 12200
rect 14424 12180 14426 12200
rect 14370 12144 14426 12180
rect 14830 12552 14886 12608
rect 14462 10512 14518 10568
rect 14830 12280 14886 12336
rect 14278 9580 14334 9616
rect 14278 9560 14280 9580
rect 14280 9560 14332 9580
rect 14332 9560 14334 9580
rect 13634 5752 13690 5808
rect 12990 5616 13046 5672
rect 13634 4936 13690 4992
rect 13174 4528 13230 4584
rect 13266 3984 13322 4040
rect 13082 3576 13138 3632
rect 12714 3068 12716 3088
rect 12716 3068 12768 3088
rect 12768 3068 12770 3088
rect 12714 3032 12770 3068
rect 13726 3848 13782 3904
rect 14370 8372 14372 8392
rect 14372 8372 14424 8392
rect 14424 8372 14426 8392
rect 14370 8336 14426 8372
rect 14646 8472 14702 8528
rect 15014 12144 15070 12200
rect 15014 11500 15016 11520
rect 15016 11500 15068 11520
rect 15068 11500 15070 11520
rect 15014 11464 15070 11500
rect 14922 10648 14978 10704
rect 14922 8916 14924 8936
rect 14924 8916 14976 8936
rect 14976 8916 14978 8936
rect 14922 8880 14978 8916
rect 14922 8744 14978 8800
rect 14830 7248 14886 7304
rect 14278 6316 14334 6352
rect 14278 6296 14280 6316
rect 14280 6296 14332 6316
rect 14332 6296 14334 6316
rect 14370 5636 14426 5672
rect 14370 5616 14372 5636
rect 14372 5616 14424 5636
rect 14424 5616 14426 5636
rect 14278 5480 14334 5536
rect 14922 5888 14978 5944
rect 16118 15544 16174 15600
rect 15198 11736 15254 11792
rect 16026 13812 16028 13832
rect 16028 13812 16080 13832
rect 16080 13812 16082 13832
rect 16026 13776 16082 13812
rect 15474 12280 15530 12336
rect 15566 11872 15622 11928
rect 15566 10668 15622 10704
rect 15566 10648 15568 10668
rect 15568 10648 15620 10668
rect 15620 10648 15622 10668
rect 15198 7284 15200 7304
rect 15200 7284 15252 7304
rect 15252 7284 15254 7304
rect 15198 7248 15254 7284
rect 15290 6840 15346 6896
rect 15658 8780 15660 8800
rect 15660 8780 15712 8800
rect 15712 8780 15714 8800
rect 15658 8744 15714 8780
rect 15750 8492 15806 8528
rect 15750 8472 15752 8492
rect 15752 8472 15804 8492
rect 15804 8472 15806 8492
rect 16118 9288 16174 9344
rect 16118 9016 16174 9072
rect 16578 10376 16634 10432
rect 16486 9560 16542 9616
rect 17222 15564 17278 15600
rect 17222 15544 17224 15564
rect 17224 15544 17276 15564
rect 17276 15544 17278 15564
rect 16762 11600 16818 11656
rect 17958 15020 18014 15056
rect 17958 15000 17960 15020
rect 17960 15000 18012 15020
rect 18012 15000 18014 15020
rect 17590 13776 17646 13832
rect 17958 14320 18014 14376
rect 18050 13640 18106 13696
rect 17222 11192 17278 11248
rect 17958 7520 18014 7576
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 9857 17778 9923 17781
rect 10501 17778 10567 17781
rect 9857 17776 10567 17778
rect 9857 17720 9862 17776
rect 9918 17720 10506 17776
rect 10562 17720 10567 17776
rect 9857 17718 10567 17720
rect 9857 17715 9923 17718
rect 10501 17715 10567 17718
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 9673 16690 9739 16693
rect 10869 16690 10935 16693
rect 12065 16690 12131 16693
rect 9673 16688 12131 16690
rect 9673 16632 9678 16688
rect 9734 16632 10874 16688
rect 10930 16632 12070 16688
rect 12126 16632 12131 16688
rect 9673 16630 12131 16632
rect 9673 16627 9739 16630
rect 10869 16627 10935 16630
rect 12065 16627 12131 16630
rect 5349 16554 5415 16557
rect 5574 16554 5580 16556
rect 5349 16552 5580 16554
rect 5349 16496 5354 16552
rect 5410 16496 5580 16552
rect 5349 16494 5580 16496
rect 5349 16491 5415 16494
rect 5574 16492 5580 16494
rect 5644 16492 5650 16556
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 8753 16282 8819 16285
rect 12617 16282 12683 16285
rect 8753 16280 12683 16282
rect 8753 16224 8758 16280
rect 8814 16224 12622 16280
rect 12678 16224 12683 16280
rect 8753 16222 12683 16224
rect 8753 16219 8819 16222
rect 12617 16219 12683 16222
rect 3049 16146 3115 16149
rect 5257 16146 5323 16149
rect 6361 16146 6427 16149
rect 9581 16146 9647 16149
rect 3049 16144 9647 16146
rect 3049 16088 3054 16144
rect 3110 16088 5262 16144
rect 5318 16088 6366 16144
rect 6422 16088 9586 16144
rect 9642 16088 9647 16144
rect 3049 16086 9647 16088
rect 3049 16083 3115 16086
rect 5257 16083 5323 16086
rect 6361 16083 6427 16086
rect 9581 16083 9647 16086
rect 9857 16146 9923 16149
rect 12893 16146 12959 16149
rect 9857 16144 12959 16146
rect 9857 16088 9862 16144
rect 9918 16088 12898 16144
rect 12954 16088 12959 16144
rect 9857 16086 12959 16088
rect 9857 16083 9923 16086
rect 12893 16083 12959 16086
rect 5073 16010 5139 16013
rect 5533 16010 5599 16013
rect 9305 16012 9371 16013
rect 5073 16008 5599 16010
rect 5073 15952 5078 16008
rect 5134 15952 5538 16008
rect 5594 15952 5599 16008
rect 5073 15950 5599 15952
rect 5073 15947 5139 15950
rect 5533 15947 5599 15950
rect 9254 15948 9260 16012
rect 9324 16010 9371 16012
rect 16481 16010 16547 16013
rect 9324 16008 16547 16010
rect 9366 15952 16486 16008
rect 16542 15952 16547 16008
rect 9324 15950 16547 15952
rect 9324 15948 9371 15950
rect 9305 15947 9371 15948
rect 16481 15947 16547 15950
rect 8937 15876 9003 15877
rect 8886 15812 8892 15876
rect 8956 15874 9003 15876
rect 9581 15874 9647 15877
rect 9949 15874 10015 15877
rect 8956 15872 9048 15874
rect 8998 15816 9048 15872
rect 8956 15814 9048 15816
rect 9581 15872 10015 15874
rect 9581 15816 9586 15872
rect 9642 15816 9954 15872
rect 10010 15816 10015 15872
rect 9581 15814 10015 15816
rect 8956 15812 9003 15814
rect 8937 15811 9003 15812
rect 9581 15811 9647 15814
rect 9949 15811 10015 15814
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 6678 15738 6684 15740
rect 4662 15678 6684 15738
rect 2957 15602 3023 15605
rect 4662 15602 4722 15678
rect 6678 15676 6684 15678
rect 6748 15738 6754 15740
rect 11329 15738 11395 15741
rect 6748 15736 11395 15738
rect 6748 15680 11334 15736
rect 11390 15680 11395 15736
rect 6748 15678 11395 15680
rect 6748 15676 6754 15678
rect 11329 15675 11395 15678
rect 2957 15600 4722 15602
rect 2957 15544 2962 15600
rect 3018 15544 4722 15600
rect 2957 15542 4722 15544
rect 7741 15602 7807 15605
rect 8569 15602 8635 15605
rect 8937 15602 9003 15605
rect 7741 15600 9003 15602
rect 7741 15544 7746 15600
rect 7802 15544 8574 15600
rect 8630 15544 8942 15600
rect 8998 15544 9003 15600
rect 7741 15542 9003 15544
rect 2957 15539 3023 15542
rect 7741 15539 7807 15542
rect 8569 15539 8635 15542
rect 8937 15539 9003 15542
rect 13445 15602 13511 15605
rect 16113 15602 16179 15605
rect 17217 15602 17283 15605
rect 13445 15600 17283 15602
rect 13445 15544 13450 15600
rect 13506 15544 16118 15600
rect 16174 15544 17222 15600
rect 17278 15544 17283 15600
rect 13445 15542 17283 15544
rect 13445 15539 13511 15542
rect 16113 15539 16179 15542
rect 17217 15539 17283 15542
rect 4613 15468 4679 15469
rect 4613 15466 4660 15468
rect 4568 15464 4660 15466
rect 4568 15408 4618 15464
rect 4568 15406 4660 15408
rect 4613 15404 4660 15406
rect 4724 15404 4730 15468
rect 5073 15466 5139 15469
rect 6085 15466 6151 15469
rect 5073 15464 6151 15466
rect 5073 15408 5078 15464
rect 5134 15408 6090 15464
rect 6146 15408 6151 15464
rect 5073 15406 6151 15408
rect 4613 15403 4679 15404
rect 5073 15403 5139 15406
rect 6085 15403 6151 15406
rect 6269 15466 6335 15469
rect 6453 15466 6519 15469
rect 7833 15466 7899 15469
rect 6269 15464 7899 15466
rect 6269 15408 6274 15464
rect 6330 15408 6458 15464
rect 6514 15408 7838 15464
rect 7894 15408 7899 15464
rect 6269 15406 7899 15408
rect 6269 15403 6335 15406
rect 6453 15403 6519 15406
rect 7833 15403 7899 15406
rect 9305 15466 9371 15469
rect 9949 15466 10015 15469
rect 9305 15464 10015 15466
rect 9305 15408 9310 15464
rect 9366 15408 9954 15464
rect 10010 15408 10015 15464
rect 9305 15406 10015 15408
rect 9305 15403 9371 15406
rect 9949 15403 10015 15406
rect 14774 15404 14780 15468
rect 14844 15466 14850 15468
rect 14917 15466 14983 15469
rect 14844 15464 14983 15466
rect 14844 15408 14922 15464
rect 14978 15408 14983 15464
rect 14844 15406 14983 15408
rect 14844 15404 14850 15406
rect 14917 15403 14983 15406
rect 8201 15330 8267 15333
rect 9581 15330 9647 15333
rect 8201 15328 9647 15330
rect 8201 15272 8206 15328
rect 8262 15272 9586 15328
rect 9642 15272 9647 15328
rect 8201 15270 9647 15272
rect 8201 15267 8267 15270
rect 9581 15267 9647 15270
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 3509 15058 3575 15061
rect 5533 15058 5599 15061
rect 3509 15056 5599 15058
rect 3509 15000 3514 15056
rect 3570 15000 5538 15056
rect 5594 15000 5599 15056
rect 3509 14998 5599 15000
rect 3509 14995 3575 14998
rect 5533 14995 5599 14998
rect 9397 15058 9463 15061
rect 9622 15058 9628 15060
rect 9397 15056 9628 15058
rect 9397 15000 9402 15056
rect 9458 15000 9628 15056
rect 9397 14998 9628 15000
rect 9397 14995 9463 14998
rect 9622 14996 9628 14998
rect 9692 14996 9698 15060
rect 10225 15058 10291 15061
rect 12801 15058 12867 15061
rect 10225 15056 12867 15058
rect 10225 15000 10230 15056
rect 10286 15000 12806 15056
rect 12862 15000 12867 15056
rect 10225 14998 12867 15000
rect 10225 14995 10291 14998
rect 12801 14995 12867 14998
rect 17953 15058 18019 15061
rect 18760 15058 19560 15088
rect 17953 15056 19560 15058
rect 17953 15000 17958 15056
rect 18014 15000 19560 15056
rect 17953 14998 19560 15000
rect 17953 14995 18019 14998
rect 18760 14968 19560 14998
rect 3233 14922 3299 14925
rect 9213 14922 9279 14925
rect 9397 14924 9463 14925
rect 9397 14922 9444 14924
rect 3233 14920 9444 14922
rect 9508 14922 9514 14924
rect 3233 14864 3238 14920
rect 3294 14864 9218 14920
rect 9274 14864 9402 14920
rect 3233 14862 9444 14864
rect 3233 14859 3299 14862
rect 9213 14859 9279 14862
rect 9397 14860 9444 14862
rect 9508 14862 9590 14922
rect 9508 14860 9514 14862
rect 9397 14859 9463 14860
rect 6821 14786 6887 14789
rect 7966 14786 7972 14788
rect 6821 14784 7972 14786
rect 6821 14728 6826 14784
rect 6882 14728 7972 14784
rect 6821 14726 7972 14728
rect 6821 14723 6887 14726
rect 7966 14724 7972 14726
rect 8036 14786 8042 14788
rect 8201 14786 8267 14789
rect 8036 14784 8267 14786
rect 8036 14728 8206 14784
rect 8262 14728 8267 14784
rect 8036 14726 8267 14728
rect 8036 14724 8042 14726
rect 8201 14723 8267 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 841 14514 907 14517
rect 798 14512 907 14514
rect 798 14456 846 14512
rect 902 14456 907 14512
rect 798 14451 907 14456
rect 9949 14514 10015 14517
rect 12341 14514 12407 14517
rect 9949 14512 12407 14514
rect 9949 14456 9954 14512
rect 10010 14456 12346 14512
rect 12402 14456 12407 14512
rect 9949 14454 12407 14456
rect 9949 14451 10015 14454
rect 12341 14451 12407 14454
rect 15101 14514 15167 14517
rect 15510 14514 15516 14516
rect 15101 14512 15516 14514
rect 15101 14456 15106 14512
rect 15162 14456 15516 14512
rect 15101 14454 15516 14456
rect 15101 14451 15167 14454
rect 15510 14452 15516 14454
rect 15580 14452 15586 14516
rect 798 14408 858 14451
rect 0 14318 858 14408
rect 0 14288 800 14318
rect 3918 14316 3924 14380
rect 3988 14378 3994 14380
rect 4705 14378 4771 14381
rect 8569 14378 8635 14381
rect 9489 14378 9555 14381
rect 3988 14376 9555 14378
rect 3988 14320 4710 14376
rect 4766 14320 8574 14376
rect 8630 14320 9494 14376
rect 9550 14320 9555 14376
rect 3988 14318 9555 14320
rect 3988 14316 3994 14318
rect 4705 14315 4771 14318
rect 8569 14315 8635 14318
rect 9489 14315 9555 14318
rect 9673 14378 9739 14381
rect 12382 14378 12388 14380
rect 9673 14376 12388 14378
rect 9673 14320 9678 14376
rect 9734 14320 12388 14376
rect 9673 14318 12388 14320
rect 9673 14315 9739 14318
rect 12382 14316 12388 14318
rect 12452 14316 12458 14380
rect 17953 14378 18019 14381
rect 18760 14378 19560 14408
rect 17953 14376 19560 14378
rect 17953 14320 17958 14376
rect 18014 14320 19560 14376
rect 17953 14318 19560 14320
rect 17953 14315 18019 14318
rect 18760 14288 19560 14318
rect 6177 14242 6243 14245
rect 6913 14242 6979 14245
rect 7046 14242 7052 14244
rect 6177 14240 7052 14242
rect 6177 14184 6182 14240
rect 6238 14184 6918 14240
rect 6974 14184 7052 14240
rect 6177 14182 7052 14184
rect 6177 14179 6243 14182
rect 6913 14179 6979 14182
rect 7046 14180 7052 14182
rect 7116 14180 7122 14244
rect 11329 14242 11395 14245
rect 13261 14242 13327 14245
rect 11329 14240 13327 14242
rect 11329 14184 11334 14240
rect 11390 14184 13266 14240
rect 13322 14184 13327 14240
rect 11329 14182 13327 14184
rect 11329 14179 11395 14182
rect 13261 14179 13327 14182
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 6126 14044 6132 14108
rect 6196 14106 6202 14108
rect 9581 14106 9647 14109
rect 6196 14104 9647 14106
rect 6196 14048 9586 14104
rect 9642 14048 9647 14104
rect 6196 14046 9647 14048
rect 6196 14044 6202 14046
rect 9581 14043 9647 14046
rect 4654 13908 4660 13972
rect 4724 13970 4730 13972
rect 5717 13970 5783 13973
rect 9857 13970 9923 13973
rect 4724 13968 5783 13970
rect 4724 13912 5722 13968
rect 5778 13912 5783 13968
rect 4724 13910 5783 13912
rect 4724 13908 4730 13910
rect 5717 13907 5783 13910
rect 5950 13968 9923 13970
rect 5950 13912 9862 13968
rect 9918 13912 9923 13968
rect 5950 13910 9923 13912
rect 4061 13834 4127 13837
rect 5950 13834 6010 13910
rect 9857 13907 9923 13910
rect 10409 13970 10475 13973
rect 10409 13968 16498 13970
rect 10409 13912 10414 13968
rect 10470 13912 16498 13968
rect 10409 13910 16498 13912
rect 10409 13907 10475 13910
rect 4061 13832 6010 13834
rect 4061 13776 4066 13832
rect 4122 13776 6010 13832
rect 4061 13774 6010 13776
rect 6177 13834 6243 13837
rect 6494 13834 6500 13836
rect 6177 13832 6500 13834
rect 6177 13776 6182 13832
rect 6238 13776 6500 13832
rect 6177 13774 6500 13776
rect 4061 13771 4127 13774
rect 6177 13771 6243 13774
rect 6494 13772 6500 13774
rect 6564 13772 6570 13836
rect 6913 13834 6979 13837
rect 9806 13834 9812 13836
rect 6913 13832 9812 13834
rect 6913 13776 6918 13832
rect 6974 13776 9812 13832
rect 6913 13774 9812 13776
rect 6913 13771 6979 13774
rect 9806 13772 9812 13774
rect 9876 13834 9882 13836
rect 10225 13834 10291 13837
rect 9876 13832 10291 13834
rect 9876 13776 10230 13832
rect 10286 13776 10291 13832
rect 9876 13774 10291 13776
rect 9876 13772 9882 13774
rect 10225 13771 10291 13774
rect 16021 13836 16087 13837
rect 16438 13836 16498 13910
rect 16021 13832 16068 13836
rect 16132 13834 16138 13836
rect 16021 13776 16026 13832
rect 16021 13772 16068 13776
rect 16132 13774 16178 13834
rect 16132 13772 16138 13774
rect 16430 13772 16436 13836
rect 16500 13834 16506 13836
rect 17585 13834 17651 13837
rect 16500 13832 17651 13834
rect 16500 13776 17590 13832
rect 17646 13776 17651 13832
rect 16500 13774 17651 13776
rect 16500 13772 16506 13774
rect 16021 13771 16087 13772
rect 17585 13771 17651 13774
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 18045 13698 18111 13701
rect 18760 13698 19560 13728
rect 18045 13696 19560 13698
rect 18045 13640 18050 13696
rect 18106 13640 19560 13696
rect 18045 13638 19560 13640
rect 18045 13635 18111 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 18760 13608 19560 13638
rect 4210 13567 4526 13568
rect 4889 13562 4955 13565
rect 7189 13562 7255 13565
rect 4889 13560 7255 13562
rect 4889 13504 4894 13560
rect 4950 13504 7194 13560
rect 7250 13504 7255 13560
rect 4889 13502 7255 13504
rect 4889 13499 4955 13502
rect 7189 13499 7255 13502
rect 9673 13562 9739 13565
rect 10409 13562 10475 13565
rect 9673 13560 10475 13562
rect 9673 13504 9678 13560
rect 9734 13504 10414 13560
rect 10470 13504 10475 13560
rect 9673 13502 10475 13504
rect 9673 13499 9739 13502
rect 10409 13499 10475 13502
rect 2497 13426 2563 13429
rect 9765 13426 9831 13429
rect 2497 13424 9831 13426
rect 2497 13368 2502 13424
rect 2558 13368 9770 13424
rect 9826 13368 9831 13424
rect 2497 13366 9831 13368
rect 2497 13363 2563 13366
rect 2730 13157 2790 13366
rect 9765 13363 9831 13366
rect 10501 13426 10567 13429
rect 14549 13426 14615 13429
rect 10501 13424 14615 13426
rect 10501 13368 10506 13424
rect 10562 13368 14554 13424
rect 14610 13368 14615 13424
rect 10501 13366 14615 13368
rect 10501 13363 10567 13366
rect 14549 13363 14615 13366
rect 2865 13290 2931 13293
rect 3141 13292 3207 13293
rect 3141 13290 3188 13292
rect 2865 13288 3188 13290
rect 2865 13232 2870 13288
rect 2926 13232 3146 13288
rect 2865 13230 3188 13232
rect 2865 13227 2931 13230
rect 3141 13228 3188 13230
rect 3252 13228 3258 13292
rect 5717 13290 5783 13293
rect 8569 13290 8635 13293
rect 5717 13288 8635 13290
rect 5717 13232 5722 13288
rect 5778 13232 8574 13288
rect 8630 13232 8635 13288
rect 5717 13230 8635 13232
rect 3141 13227 3207 13228
rect 5717 13227 5783 13230
rect 8569 13227 8635 13230
rect 12566 13228 12572 13292
rect 12636 13290 12642 13292
rect 12985 13290 13051 13293
rect 12636 13288 13051 13290
rect 12636 13232 12990 13288
rect 13046 13232 13051 13288
rect 12636 13230 13051 13232
rect 12636 13228 12642 13230
rect 12985 13227 13051 13230
rect 2730 13152 2839 13157
rect 11329 13156 11395 13157
rect 11278 13154 11284 13156
rect 2730 13096 2778 13152
rect 2834 13096 2839 13152
rect 2730 13094 2839 13096
rect 11238 13094 11284 13154
rect 11348 13152 11395 13156
rect 11390 13096 11395 13152
rect 2773 13091 2839 13094
rect 11278 13092 11284 13094
rect 11348 13092 11395 13096
rect 11329 13091 11395 13092
rect 11513 13154 11579 13157
rect 11646 13154 11652 13156
rect 11513 13152 11652 13154
rect 11513 13096 11518 13152
rect 11574 13096 11652 13152
rect 11513 13094 11652 13096
rect 11513 13091 11579 13094
rect 11646 13092 11652 13094
rect 11716 13092 11722 13156
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 9765 13018 9831 13021
rect 12341 13018 12407 13021
rect 9765 13016 12407 13018
rect 9765 12960 9770 13016
rect 9826 12960 12346 13016
rect 12402 12960 12407 13016
rect 9765 12958 12407 12960
rect 9765 12955 9831 12958
rect 12341 12955 12407 12958
rect 5993 12882 6059 12885
rect 11881 12882 11947 12885
rect 5993 12880 14060 12882
rect 5993 12824 5998 12880
rect 6054 12824 11886 12880
rect 11942 12824 14060 12880
rect 5993 12822 14060 12824
rect 5993 12819 6059 12822
rect 11881 12819 11947 12822
rect 4889 12746 4955 12749
rect 5758 12746 5764 12748
rect 4889 12744 5764 12746
rect 4889 12688 4894 12744
rect 4950 12688 5764 12744
rect 4889 12686 5764 12688
rect 4889 12683 4955 12686
rect 5758 12684 5764 12686
rect 5828 12684 5834 12748
rect 6913 12746 6979 12749
rect 7414 12746 7420 12748
rect 6913 12744 7420 12746
rect 6913 12688 6918 12744
rect 6974 12688 7420 12744
rect 6913 12686 7420 12688
rect 3049 12612 3115 12613
rect 2998 12610 3004 12612
rect 2958 12550 3004 12610
rect 3068 12608 3115 12612
rect 3110 12552 3115 12608
rect 2998 12548 3004 12550
rect 3068 12548 3115 12552
rect 5766 12610 5826 12684
rect 6913 12683 6979 12686
rect 7414 12684 7420 12686
rect 7484 12684 7490 12748
rect 10685 12746 10751 12749
rect 13353 12746 13419 12749
rect 10685 12744 13419 12746
rect 10685 12688 10690 12744
rect 10746 12688 13358 12744
rect 13414 12688 13419 12744
rect 10685 12686 13419 12688
rect 14000 12746 14060 12822
rect 14457 12746 14523 12749
rect 15142 12746 15148 12748
rect 14000 12744 15148 12746
rect 14000 12688 14462 12744
rect 14518 12688 15148 12744
rect 14000 12686 15148 12688
rect 10685 12683 10751 12686
rect 13353 12683 13419 12686
rect 14457 12683 14523 12686
rect 15142 12684 15148 12686
rect 15212 12684 15218 12748
rect 7741 12610 7807 12613
rect 5766 12608 7807 12610
rect 5766 12552 7746 12608
rect 7802 12552 7807 12608
rect 5766 12550 7807 12552
rect 3049 12547 3115 12548
rect 7741 12547 7807 12550
rect 11605 12610 11671 12613
rect 14089 12610 14155 12613
rect 14825 12610 14891 12613
rect 11605 12608 14891 12610
rect 11605 12552 11610 12608
rect 11666 12552 14094 12608
rect 14150 12552 14830 12608
rect 14886 12552 14891 12608
rect 11605 12550 14891 12552
rect 11605 12547 11671 12550
rect 14089 12547 14155 12550
rect 14825 12547 14891 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 5073 12474 5139 12477
rect 7230 12474 7236 12476
rect 5073 12472 7236 12474
rect 5073 12416 5078 12472
rect 5134 12416 7236 12472
rect 5073 12414 7236 12416
rect 5073 12411 5139 12414
rect 7230 12412 7236 12414
rect 7300 12412 7306 12476
rect 9070 12412 9076 12476
rect 9140 12474 9146 12476
rect 9489 12474 9555 12477
rect 9140 12472 9555 12474
rect 9140 12416 9494 12472
rect 9550 12416 9555 12472
rect 9140 12414 9555 12416
rect 9140 12412 9146 12414
rect 9489 12411 9555 12414
rect 9765 12474 9831 12477
rect 10777 12474 10843 12477
rect 9765 12472 10843 12474
rect 9765 12416 9770 12472
rect 9826 12416 10782 12472
rect 10838 12416 10843 12472
rect 9765 12414 10843 12416
rect 9765 12411 9831 12414
rect 10777 12411 10843 12414
rect 11237 12474 11303 12477
rect 13353 12474 13419 12477
rect 11237 12472 13419 12474
rect 11237 12416 11242 12472
rect 11298 12416 13358 12472
rect 13414 12416 13419 12472
rect 11237 12414 13419 12416
rect 11237 12411 11303 12414
rect 13353 12411 13419 12414
rect 8569 12338 8635 12341
rect 11697 12338 11763 12341
rect 14825 12338 14891 12341
rect 15469 12338 15535 12341
rect 8569 12336 15535 12338
rect 8569 12280 8574 12336
rect 8630 12280 11702 12336
rect 11758 12280 14830 12336
rect 14886 12280 15474 12336
rect 15530 12280 15535 12336
rect 8569 12278 15535 12280
rect 8569 12275 8635 12278
rect 11697 12275 11763 12278
rect 14825 12275 14891 12278
rect 15469 12275 15535 12278
rect 4521 12202 4587 12205
rect 5390 12202 5396 12204
rect 4521 12200 5396 12202
rect 4521 12144 4526 12200
rect 4582 12144 5396 12200
rect 4521 12142 5396 12144
rect 4521 12139 4587 12142
rect 5390 12140 5396 12142
rect 5460 12202 5466 12204
rect 12525 12202 12591 12205
rect 14365 12204 14431 12205
rect 15009 12204 15075 12205
rect 14365 12202 14412 12204
rect 5460 12200 12591 12202
rect 5460 12144 12530 12200
rect 12586 12144 12591 12200
rect 5460 12142 12591 12144
rect 14320 12200 14412 12202
rect 14320 12144 14370 12200
rect 14320 12142 14412 12144
rect 5460 12140 5466 12142
rect 12525 12139 12591 12142
rect 14365 12140 14412 12142
rect 14476 12140 14482 12204
rect 14958 12140 14964 12204
rect 15028 12202 15075 12204
rect 15028 12200 15120 12202
rect 15070 12144 15120 12200
rect 15028 12142 15120 12144
rect 15028 12140 15075 12142
rect 14365 12139 14431 12140
rect 15009 12139 15075 12140
rect 8569 12066 8635 12069
rect 8937 12066 9003 12069
rect 8569 12064 9003 12066
rect 8569 12008 8574 12064
rect 8630 12008 8942 12064
rect 8998 12008 9003 12064
rect 8569 12006 9003 12008
rect 8569 12003 8635 12006
rect 8937 12003 9003 12006
rect 9765 12066 9831 12069
rect 12985 12066 13051 12069
rect 9765 12064 13051 12066
rect 9765 12008 9770 12064
rect 9826 12008 12990 12064
rect 13046 12008 13051 12064
rect 9765 12006 13051 12008
rect 9765 12003 9831 12006
rect 12985 12003 13051 12006
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 8334 11868 8340 11932
rect 8404 11930 8410 11932
rect 11053 11930 11119 11933
rect 8404 11928 11119 11930
rect 8404 11872 11058 11928
rect 11114 11872 11119 11928
rect 8404 11870 11119 11872
rect 8404 11868 8410 11870
rect 11053 11867 11119 11870
rect 12249 11930 12315 11933
rect 15561 11930 15627 11933
rect 12249 11928 15627 11930
rect 12249 11872 12254 11928
rect 12310 11872 15566 11928
rect 15622 11872 15627 11928
rect 12249 11870 15627 11872
rect 12249 11867 12315 11870
rect 15561 11867 15627 11870
rect 5073 11794 5139 11797
rect 15193 11794 15259 11797
rect 15326 11794 15332 11796
rect 5073 11792 15332 11794
rect 5073 11736 5078 11792
rect 5134 11736 15198 11792
rect 15254 11736 15332 11792
rect 5073 11734 15332 11736
rect 5073 11731 5139 11734
rect 15193 11731 15259 11734
rect 15326 11732 15332 11734
rect 15396 11732 15402 11796
rect 8293 11658 8359 11661
rect 9857 11658 9923 11661
rect 8293 11656 9923 11658
rect 8293 11600 8298 11656
rect 8354 11600 9862 11656
rect 9918 11600 9923 11656
rect 8293 11598 9923 11600
rect 8293 11595 8359 11598
rect 9857 11595 9923 11598
rect 10041 11658 10107 11661
rect 12433 11658 12499 11661
rect 16757 11658 16823 11661
rect 10041 11656 16823 11658
rect 10041 11600 10046 11656
rect 10102 11600 12438 11656
rect 12494 11600 16762 11656
rect 16818 11600 16823 11656
rect 10041 11598 16823 11600
rect 10041 11595 10107 11598
rect 12433 11595 12499 11598
rect 16757 11595 16823 11598
rect 7925 11522 7991 11525
rect 9581 11522 9647 11525
rect 7925 11520 9647 11522
rect 7925 11464 7930 11520
rect 7986 11464 9586 11520
rect 9642 11464 9647 11520
rect 7925 11462 9647 11464
rect 7925 11459 7991 11462
rect 9581 11459 9647 11462
rect 9765 11522 9831 11525
rect 10225 11522 10291 11525
rect 9765 11520 10291 11522
rect 9765 11464 9770 11520
rect 9826 11464 10230 11520
rect 10286 11464 10291 11520
rect 9765 11462 10291 11464
rect 9765 11459 9831 11462
rect 10225 11459 10291 11462
rect 13721 11522 13787 11525
rect 15009 11522 15075 11525
rect 13721 11520 15075 11522
rect 13721 11464 13726 11520
rect 13782 11464 15014 11520
rect 15070 11464 15075 11520
rect 13721 11462 15075 11464
rect 13721 11459 13787 11462
rect 15009 11459 15075 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 9673 11386 9739 11389
rect 10317 11386 10383 11389
rect 9673 11384 10383 11386
rect 9673 11328 9678 11384
rect 9734 11328 10322 11384
rect 10378 11328 10383 11384
rect 9673 11326 10383 11328
rect 9673 11323 9739 11326
rect 10317 11323 10383 11326
rect 10501 11386 10567 11389
rect 12893 11386 12959 11389
rect 10501 11384 12959 11386
rect 10501 11328 10506 11384
rect 10562 11328 12898 11384
rect 12954 11328 12959 11384
rect 10501 11326 12959 11328
rect 10501 11323 10567 11326
rect 12893 11323 12959 11326
rect 6913 11252 6979 11253
rect 6862 11250 6868 11252
rect 6822 11190 6868 11250
rect 6932 11248 6979 11252
rect 6974 11192 6979 11248
rect 6862 11188 6868 11190
rect 6932 11188 6979 11192
rect 6913 11187 6979 11188
rect 9121 11250 9187 11253
rect 11278 11250 11284 11252
rect 9121 11248 11284 11250
rect 9121 11192 9126 11248
rect 9182 11192 11284 11248
rect 9121 11190 11284 11192
rect 9121 11187 9187 11190
rect 11278 11188 11284 11190
rect 11348 11250 11354 11252
rect 17217 11250 17283 11253
rect 11348 11248 17283 11250
rect 11348 11192 17222 11248
rect 17278 11192 17283 11248
rect 11348 11190 17283 11192
rect 11348 11188 11354 11190
rect 17217 11187 17283 11190
rect 2589 11114 2655 11117
rect 6085 11114 6151 11117
rect 2589 11112 6151 11114
rect 2589 11056 2594 11112
rect 2650 11056 6090 11112
rect 6146 11056 6151 11112
rect 2589 11054 6151 11056
rect 2589 11051 2655 11054
rect 6085 11051 6151 11054
rect 6678 11052 6684 11116
rect 6748 11114 6754 11116
rect 6821 11114 6887 11117
rect 10910 11114 10916 11116
rect 6748 11112 10916 11114
rect 6748 11056 6826 11112
rect 6882 11056 10916 11112
rect 6748 11054 10916 11056
rect 6748 11052 6754 11054
rect 6821 11051 6887 11054
rect 10910 11052 10916 11054
rect 10980 11114 10986 11116
rect 12065 11114 12131 11117
rect 10980 11112 12131 11114
rect 10980 11056 12070 11112
rect 12126 11056 12131 11112
rect 10980 11054 12131 11056
rect 10980 11052 10986 11054
rect 12065 11051 12131 11054
rect 12801 11114 12867 11117
rect 13302 11114 13308 11116
rect 12801 11112 13308 11114
rect 12801 11056 12806 11112
rect 12862 11056 13308 11112
rect 12801 11054 13308 11056
rect 12801 11051 12867 11054
rect 13302 11052 13308 11054
rect 13372 11052 13378 11116
rect 8334 10916 8340 10980
rect 8404 10978 8410 10980
rect 8753 10978 8819 10981
rect 8404 10976 8819 10978
rect 8404 10920 8758 10976
rect 8814 10920 8819 10976
rect 8404 10918 8819 10920
rect 8404 10916 8410 10918
rect 8753 10915 8819 10918
rect 11646 10916 11652 10980
rect 11716 10978 11722 10980
rect 12525 10978 12591 10981
rect 11716 10976 12591 10978
rect 11716 10920 12530 10976
rect 12586 10920 12591 10976
rect 11716 10918 12591 10920
rect 11716 10916 11722 10918
rect 12525 10915 12591 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 6494 10780 6500 10844
rect 6564 10842 6570 10844
rect 11881 10842 11947 10845
rect 6564 10840 11947 10842
rect 6564 10784 11886 10840
rect 11942 10784 11947 10840
rect 6564 10782 11947 10784
rect 6564 10780 6570 10782
rect 11881 10779 11947 10782
rect 8753 10706 8819 10709
rect 9213 10706 9279 10709
rect 8753 10704 9279 10706
rect 8753 10648 8758 10704
rect 8814 10648 9218 10704
rect 9274 10648 9279 10704
rect 8753 10646 9279 10648
rect 8753 10643 8819 10646
rect 9213 10643 9279 10646
rect 10133 10706 10199 10709
rect 11053 10706 11119 10709
rect 12985 10706 13051 10709
rect 10133 10704 13051 10706
rect 10133 10648 10138 10704
rect 10194 10648 11058 10704
rect 11114 10648 12990 10704
rect 13046 10648 13051 10704
rect 10133 10646 13051 10648
rect 10133 10643 10199 10646
rect 11053 10643 11119 10646
rect 12985 10643 13051 10646
rect 13261 10706 13327 10709
rect 13486 10706 13492 10708
rect 13261 10704 13492 10706
rect 13261 10648 13266 10704
rect 13322 10648 13492 10704
rect 13261 10646 13492 10648
rect 13261 10643 13327 10646
rect 13486 10644 13492 10646
rect 13556 10706 13562 10708
rect 13997 10706 14063 10709
rect 14917 10708 14983 10709
rect 14917 10706 14964 10708
rect 13556 10704 14063 10706
rect 13556 10648 14002 10704
rect 14058 10648 14063 10704
rect 13556 10646 14063 10648
rect 14872 10704 14964 10706
rect 14872 10648 14922 10704
rect 14872 10646 14964 10648
rect 13556 10644 13562 10646
rect 13997 10643 14063 10646
rect 14917 10644 14964 10646
rect 15028 10644 15034 10708
rect 15142 10644 15148 10708
rect 15212 10706 15218 10708
rect 15561 10706 15627 10709
rect 15212 10704 15627 10706
rect 15212 10648 15566 10704
rect 15622 10648 15627 10704
rect 15212 10646 15627 10648
rect 15212 10644 15218 10646
rect 14917 10643 14983 10644
rect 15561 10643 15627 10646
rect 4061 10570 4127 10573
rect 4654 10570 4660 10572
rect 4061 10568 4660 10570
rect 4061 10512 4066 10568
rect 4122 10512 4660 10568
rect 4061 10510 4660 10512
rect 4061 10507 4127 10510
rect 4654 10508 4660 10510
rect 4724 10508 4730 10572
rect 4981 10570 5047 10573
rect 5901 10570 5967 10573
rect 8293 10570 8359 10573
rect 11789 10570 11855 10573
rect 4981 10568 8359 10570
rect 4981 10512 4986 10568
rect 5042 10512 5906 10568
rect 5962 10512 8298 10568
rect 8354 10512 8359 10568
rect 4981 10510 8359 10512
rect 4981 10507 5047 10510
rect 5901 10507 5967 10510
rect 8293 10507 8359 10510
rect 11654 10568 11855 10570
rect 11654 10512 11794 10568
rect 11850 10512 11855 10568
rect 11654 10510 11855 10512
rect 5809 10434 5875 10437
rect 7097 10434 7163 10437
rect 5809 10432 7163 10434
rect 5809 10376 5814 10432
rect 5870 10376 7102 10432
rect 7158 10376 7163 10432
rect 5809 10374 7163 10376
rect 5809 10371 5875 10374
rect 7097 10371 7163 10374
rect 8661 10434 8727 10437
rect 11329 10434 11395 10437
rect 8661 10432 11395 10434
rect 8661 10376 8666 10432
rect 8722 10376 11334 10432
rect 11390 10376 11395 10432
rect 8661 10374 11395 10376
rect 8661 10371 8727 10374
rect 11329 10371 11395 10374
rect 11513 10434 11579 10437
rect 11654 10434 11714 10510
rect 11789 10507 11855 10510
rect 12382 10508 12388 10572
rect 12452 10570 12458 10572
rect 12709 10570 12775 10573
rect 14457 10570 14523 10573
rect 12452 10568 14523 10570
rect 12452 10512 12714 10568
rect 12770 10512 14462 10568
rect 14518 10512 14523 10568
rect 12452 10510 14523 10512
rect 12452 10508 12458 10510
rect 12709 10507 12775 10510
rect 14457 10507 14523 10510
rect 11513 10432 11714 10434
rect 11513 10376 11518 10432
rect 11574 10376 11714 10432
rect 11513 10374 11714 10376
rect 13077 10434 13143 10437
rect 16573 10434 16639 10437
rect 13077 10432 16639 10434
rect 13077 10376 13082 10432
rect 13138 10376 16578 10432
rect 16634 10376 16639 10432
rect 13077 10374 16639 10376
rect 11513 10371 11579 10374
rect 13077 10371 13143 10374
rect 16573 10371 16639 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 9070 10236 9076 10300
rect 9140 10298 9146 10300
rect 9489 10298 9555 10301
rect 9140 10296 9555 10298
rect 9140 10240 9494 10296
rect 9550 10240 9555 10296
rect 9140 10238 9555 10240
rect 9140 10236 9146 10238
rect 9489 10235 9555 10238
rect 11145 10298 11211 10301
rect 13169 10298 13235 10301
rect 11145 10296 13235 10298
rect 11145 10240 11150 10296
rect 11206 10240 13174 10296
rect 13230 10240 13235 10296
rect 11145 10238 13235 10240
rect 11145 10235 11211 10238
rect 13169 10235 13235 10238
rect 3877 10162 3943 10165
rect 4429 10162 4495 10165
rect 3877 10160 4495 10162
rect 3877 10104 3882 10160
rect 3938 10104 4434 10160
rect 4490 10104 4495 10160
rect 3877 10102 4495 10104
rect 3877 10099 3943 10102
rect 4429 10099 4495 10102
rect 10869 10162 10935 10165
rect 12433 10162 12499 10165
rect 10869 10160 12499 10162
rect 10869 10104 10874 10160
rect 10930 10104 12438 10160
rect 12494 10104 12499 10160
rect 10869 10102 12499 10104
rect 10869 10099 10935 10102
rect 12433 10099 12499 10102
rect 3918 9964 3924 10028
rect 3988 10026 3994 10028
rect 4705 10026 4771 10029
rect 3988 10024 4771 10026
rect 3988 9968 4710 10024
rect 4766 9968 4771 10024
rect 3988 9966 4771 9968
rect 3988 9964 3994 9966
rect 4705 9963 4771 9966
rect 5257 10024 5323 10029
rect 5257 9968 5262 10024
rect 5318 9968 5323 10024
rect 5257 9963 5323 9968
rect 8569 10026 8635 10029
rect 9489 10026 9555 10029
rect 8569 10024 9555 10026
rect 8569 9968 8574 10024
rect 8630 9968 9494 10024
rect 9550 9968 9555 10024
rect 8569 9966 9555 9968
rect 8569 9963 8635 9966
rect 9489 9963 9555 9966
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 3325 9756 3391 9757
rect 3325 9752 3372 9756
rect 3436 9754 3442 9756
rect 3325 9696 3330 9752
rect 3325 9692 3372 9696
rect 3436 9694 3482 9754
rect 3436 9692 3442 9694
rect 5260 9693 5320 9963
rect 5717 9890 5783 9893
rect 8569 9890 8635 9893
rect 9397 9890 9463 9893
rect 5717 9888 9463 9890
rect 5717 9832 5722 9888
rect 5778 9832 8574 9888
rect 8630 9832 9402 9888
rect 9458 9832 9463 9888
rect 5717 9830 9463 9832
rect 5717 9827 5783 9830
rect 8569 9827 8635 9830
rect 9397 9827 9463 9830
rect 7557 9754 7623 9757
rect 10593 9754 10659 9757
rect 7557 9752 10659 9754
rect 7557 9696 7562 9752
rect 7618 9696 10598 9752
rect 10654 9696 10659 9752
rect 7557 9694 10659 9696
rect 3325 9691 3391 9692
rect 5257 9688 5323 9693
rect 7557 9691 7623 9694
rect 10593 9691 10659 9694
rect 11881 9754 11947 9757
rect 12014 9754 12020 9756
rect 11881 9752 12020 9754
rect 11881 9696 11886 9752
rect 11942 9696 12020 9752
rect 11881 9694 12020 9696
rect 11881 9691 11947 9694
rect 12014 9692 12020 9694
rect 12084 9692 12090 9756
rect 5257 9632 5262 9688
rect 5318 9632 5323 9688
rect 5257 9627 5323 9632
rect 3049 9620 3115 9621
rect 2998 9556 3004 9620
rect 3068 9618 3115 9620
rect 5901 9618 5967 9621
rect 6126 9618 6132 9620
rect 3068 9616 3160 9618
rect 3110 9560 3160 9616
rect 3068 9558 3160 9560
rect 5901 9616 6132 9618
rect 5901 9560 5906 9616
rect 5962 9560 6132 9616
rect 5901 9558 6132 9560
rect 3068 9556 3115 9558
rect 3049 9555 3115 9556
rect 5901 9555 5967 9558
rect 6126 9556 6132 9558
rect 6196 9556 6202 9620
rect 6453 9618 6519 9621
rect 6637 9618 6703 9621
rect 6453 9616 6703 9618
rect 6453 9560 6458 9616
rect 6514 9560 6642 9616
rect 6698 9560 6703 9616
rect 6453 9558 6703 9560
rect 6453 9555 6519 9558
rect 6637 9555 6703 9558
rect 7230 9556 7236 9620
rect 7300 9618 7306 9620
rect 12709 9618 12775 9621
rect 7300 9616 12775 9618
rect 7300 9560 12714 9616
rect 12770 9560 12775 9616
rect 7300 9558 12775 9560
rect 7300 9556 7306 9558
rect 12709 9555 12775 9558
rect 14273 9618 14339 9621
rect 16481 9620 16547 9621
rect 14406 9618 14412 9620
rect 14273 9616 14412 9618
rect 14273 9560 14278 9616
rect 14334 9560 14412 9616
rect 14273 9558 14412 9560
rect 14273 9555 14339 9558
rect 14406 9556 14412 9558
rect 14476 9556 14482 9620
rect 16430 9618 16436 9620
rect 16390 9558 16436 9618
rect 16500 9616 16547 9620
rect 16542 9560 16547 9616
rect 16430 9556 16436 9558
rect 16500 9556 16547 9560
rect 16481 9555 16547 9556
rect 5574 9420 5580 9484
rect 5644 9482 5650 9484
rect 5809 9482 5875 9485
rect 5644 9480 5875 9482
rect 5644 9424 5814 9480
rect 5870 9424 5875 9480
rect 5644 9422 5875 9424
rect 5644 9420 5650 9422
rect 5809 9419 5875 9422
rect 9622 9420 9628 9484
rect 9692 9482 9698 9484
rect 14222 9482 14228 9484
rect 9692 9422 14228 9482
rect 9692 9420 9698 9422
rect 14222 9420 14228 9422
rect 14292 9420 14298 9484
rect 10409 9346 10475 9349
rect 12249 9346 12315 9349
rect 12433 9346 12499 9349
rect 10409 9344 12499 9346
rect 10409 9288 10414 9344
rect 10470 9288 12254 9344
rect 12310 9288 12438 9344
rect 12494 9288 12499 9344
rect 10409 9286 12499 9288
rect 10409 9283 10475 9286
rect 12249 9283 12315 9286
rect 12433 9283 12499 9286
rect 13353 9346 13419 9349
rect 16113 9348 16179 9349
rect 16062 9346 16068 9348
rect 13353 9344 16068 9346
rect 16132 9344 16179 9348
rect 13353 9288 13358 9344
rect 13414 9288 16068 9344
rect 16174 9288 16179 9344
rect 13353 9286 16068 9288
rect 13353 9283 13419 9286
rect 16062 9284 16068 9286
rect 16132 9284 16179 9288
rect 16113 9283 16179 9284
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 2957 9074 3023 9077
rect 4429 9074 4495 9077
rect 2957 9072 4495 9074
rect 2957 9016 2962 9072
rect 3018 9016 4434 9072
rect 4490 9016 4495 9072
rect 2957 9014 4495 9016
rect 2957 9011 3023 9014
rect 4429 9011 4495 9014
rect 6913 9074 6979 9077
rect 7046 9074 7052 9076
rect 6913 9072 7052 9074
rect 6913 9016 6918 9072
rect 6974 9016 7052 9072
rect 6913 9014 7052 9016
rect 6913 9011 6979 9014
rect 7046 9012 7052 9014
rect 7116 9012 7122 9076
rect 8109 9074 8175 9077
rect 11513 9074 11579 9077
rect 8109 9072 11579 9074
rect 8109 9016 8114 9072
rect 8170 9016 11518 9072
rect 11574 9016 11579 9072
rect 8109 9014 11579 9016
rect 8109 9011 8175 9014
rect 11513 9011 11579 9014
rect 12249 9074 12315 9077
rect 16113 9074 16179 9077
rect 12249 9072 16179 9074
rect 12249 9016 12254 9072
rect 12310 9016 16118 9072
rect 16174 9016 16179 9072
rect 12249 9014 16179 9016
rect 12249 9011 12315 9014
rect 16113 9011 16179 9014
rect 0 8938 800 8968
rect 1025 8938 1091 8941
rect 0 8936 1091 8938
rect 0 8880 1030 8936
rect 1086 8880 1091 8936
rect 0 8878 1091 8880
rect 0 8848 800 8878
rect 1025 8875 1091 8878
rect 2998 8876 3004 8940
rect 3068 8938 3074 8940
rect 4153 8938 4219 8941
rect 6678 8938 6684 8940
rect 3068 8936 4219 8938
rect 3068 8880 4158 8936
rect 4214 8880 4219 8936
rect 3068 8878 4219 8880
rect 3068 8876 3074 8878
rect 2773 8802 2839 8805
rect 3006 8802 3066 8876
rect 4153 8875 4219 8878
rect 4662 8878 6684 8938
rect 2773 8800 3066 8802
rect 2773 8744 2778 8800
rect 2834 8744 3066 8800
rect 2773 8742 3066 8744
rect 3785 8802 3851 8805
rect 4662 8802 4722 8878
rect 6678 8876 6684 8878
rect 6748 8876 6754 8940
rect 14774 8876 14780 8940
rect 14844 8938 14850 8940
rect 14917 8938 14983 8941
rect 14844 8936 14983 8938
rect 14844 8880 14922 8936
rect 14978 8880 14983 8936
rect 14844 8878 14983 8880
rect 14844 8876 14850 8878
rect 14917 8875 14983 8878
rect 3785 8800 4722 8802
rect 3785 8744 3790 8800
rect 3846 8744 4722 8800
rect 3785 8742 4722 8744
rect 6913 8802 6979 8805
rect 7230 8802 7236 8804
rect 6913 8800 7236 8802
rect 6913 8744 6918 8800
rect 6974 8744 7236 8800
rect 6913 8742 7236 8744
rect 2773 8739 2839 8742
rect 3785 8739 3851 8742
rect 6913 8739 6979 8742
rect 7230 8740 7236 8742
rect 7300 8740 7306 8804
rect 14917 8802 14983 8805
rect 15653 8802 15719 8805
rect 14917 8800 15719 8802
rect 14917 8744 14922 8800
rect 14978 8744 15658 8800
rect 15714 8744 15719 8800
rect 14917 8742 15719 8744
rect 14917 8739 14983 8742
rect 15653 8739 15719 8742
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 8477 8666 8543 8669
rect 10869 8666 10935 8669
rect 11881 8666 11947 8669
rect 5582 8664 11947 8666
rect 5582 8608 8482 8664
rect 8538 8608 10874 8664
rect 10930 8608 11886 8664
rect 11942 8608 11947 8664
rect 5582 8606 11947 8608
rect 3141 8530 3207 8533
rect 3785 8530 3851 8533
rect 5165 8530 5231 8533
rect 5582 8530 5642 8606
rect 8477 8603 8543 8606
rect 10869 8603 10935 8606
rect 11881 8603 11947 8606
rect 3141 8528 5642 8530
rect 3141 8472 3146 8528
rect 3202 8472 3790 8528
rect 3846 8472 5170 8528
rect 5226 8472 5642 8528
rect 3141 8470 5642 8472
rect 5993 8530 6059 8533
rect 6637 8530 6703 8533
rect 14641 8530 14707 8533
rect 5993 8528 14707 8530
rect 5993 8472 5998 8528
rect 6054 8472 6642 8528
rect 6698 8472 14646 8528
rect 14702 8472 14707 8528
rect 5993 8470 14707 8472
rect 3141 8467 3207 8470
rect 3785 8467 3851 8470
rect 5165 8467 5231 8470
rect 5993 8467 6059 8470
rect 6637 8467 6703 8470
rect 14641 8467 14707 8470
rect 15510 8468 15516 8532
rect 15580 8530 15586 8532
rect 15745 8530 15811 8533
rect 15580 8528 15811 8530
rect 15580 8472 15750 8528
rect 15806 8472 15811 8528
rect 15580 8470 15811 8472
rect 15580 8468 15586 8470
rect 15745 8467 15811 8470
rect 7189 8394 7255 8397
rect 7649 8394 7715 8397
rect 7189 8392 7715 8394
rect 7189 8336 7194 8392
rect 7250 8336 7654 8392
rect 7710 8336 7715 8392
rect 7189 8334 7715 8336
rect 7189 8331 7255 8334
rect 7649 8331 7715 8334
rect 8293 8394 8359 8397
rect 9029 8394 9095 8397
rect 9949 8394 10015 8397
rect 13670 8394 13676 8396
rect 8293 8392 10015 8394
rect 8293 8336 8298 8392
rect 8354 8336 9034 8392
rect 9090 8336 9954 8392
rect 10010 8336 10015 8392
rect 8293 8334 10015 8336
rect 8293 8331 8359 8334
rect 9029 8331 9095 8334
rect 9949 8331 10015 8334
rect 12390 8334 13676 8394
rect 7281 8258 7347 8261
rect 9254 8258 9260 8260
rect 7281 8256 9260 8258
rect 7281 8200 7286 8256
rect 7342 8200 9260 8256
rect 7281 8198 9260 8200
rect 7281 8195 7347 8198
rect 9254 8196 9260 8198
rect 9324 8196 9330 8260
rect 9806 8196 9812 8260
rect 9876 8258 9882 8260
rect 10225 8258 10291 8261
rect 12390 8258 12450 8334
rect 13670 8332 13676 8334
rect 13740 8394 13746 8396
rect 14365 8394 14431 8397
rect 13740 8392 14431 8394
rect 13740 8336 14370 8392
rect 14426 8336 14431 8392
rect 13740 8334 14431 8336
rect 13740 8332 13746 8334
rect 14365 8331 14431 8334
rect 9876 8256 12450 8258
rect 9876 8200 10230 8256
rect 10286 8200 12450 8256
rect 9876 8198 12450 8200
rect 9876 8196 9882 8198
rect 10225 8195 10291 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 6545 7986 6611 7989
rect 7649 7986 7715 7989
rect 6545 7984 7715 7986
rect 6545 7928 6550 7984
rect 6606 7928 7654 7984
rect 7710 7928 7715 7984
rect 6545 7926 7715 7928
rect 6545 7923 6611 7926
rect 7649 7923 7715 7926
rect 9213 7986 9279 7989
rect 9438 7986 9444 7988
rect 9213 7984 9444 7986
rect 9213 7928 9218 7984
rect 9274 7928 9444 7984
rect 9213 7926 9444 7928
rect 9213 7923 9279 7926
rect 9438 7924 9444 7926
rect 9508 7924 9514 7988
rect 11513 7986 11579 7989
rect 13997 7986 14063 7989
rect 11513 7984 14063 7986
rect 11513 7928 11518 7984
rect 11574 7928 14002 7984
rect 14058 7928 14063 7984
rect 11513 7926 14063 7928
rect 11513 7923 11579 7926
rect 13997 7923 14063 7926
rect 5993 7850 6059 7853
rect 8569 7850 8635 7853
rect 5993 7848 8635 7850
rect 5993 7792 5998 7848
rect 6054 7792 8574 7848
rect 8630 7792 8635 7848
rect 5993 7790 8635 7792
rect 5993 7787 6059 7790
rect 8569 7787 8635 7790
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 10685 7578 10751 7581
rect 12525 7578 12591 7581
rect 10685 7576 12591 7578
rect 10685 7520 10690 7576
rect 10746 7520 12530 7576
rect 12586 7520 12591 7576
rect 10685 7518 12591 7520
rect 10685 7515 10751 7518
rect 12525 7515 12591 7518
rect 17953 7578 18019 7581
rect 18760 7578 19560 7608
rect 17953 7576 19560 7578
rect 17953 7520 17958 7576
rect 18014 7520 19560 7576
rect 17953 7518 19560 7520
rect 17953 7515 18019 7518
rect 18760 7488 19560 7518
rect 10041 7442 10107 7445
rect 10910 7442 10916 7444
rect 10041 7440 10916 7442
rect 10041 7384 10046 7440
rect 10102 7384 10916 7440
rect 10041 7382 10916 7384
rect 10041 7379 10107 7382
rect 10910 7380 10916 7382
rect 10980 7442 10986 7444
rect 12617 7442 12683 7445
rect 10980 7440 12683 7442
rect 10980 7384 12622 7440
rect 12678 7384 12683 7440
rect 10980 7382 12683 7384
rect 10980 7380 10986 7382
rect 12617 7379 12683 7382
rect 5349 7308 5415 7309
rect 5349 7306 5396 7308
rect 5304 7304 5396 7306
rect 5304 7248 5354 7304
rect 5304 7246 5396 7248
rect 5349 7244 5396 7246
rect 5460 7244 5466 7308
rect 10174 7244 10180 7308
rect 10244 7306 10250 7308
rect 10317 7306 10383 7309
rect 10244 7304 10383 7306
rect 10244 7248 10322 7304
rect 10378 7248 10383 7304
rect 10244 7246 10383 7248
rect 10244 7244 10250 7246
rect 5349 7243 5415 7244
rect 10317 7243 10383 7246
rect 11513 7306 11579 7309
rect 14825 7306 14891 7309
rect 15193 7306 15259 7309
rect 11513 7304 15259 7306
rect 11513 7248 11518 7304
rect 11574 7248 14830 7304
rect 14886 7248 15198 7304
rect 15254 7248 15259 7304
rect 11513 7246 15259 7248
rect 11513 7243 11579 7246
rect 14825 7243 14891 7246
rect 15193 7243 15259 7246
rect 10961 7170 11027 7173
rect 12801 7170 12867 7173
rect 13261 7170 13327 7173
rect 10961 7168 13327 7170
rect 10961 7112 10966 7168
rect 11022 7112 12806 7168
rect 12862 7112 13266 7168
rect 13322 7112 13327 7168
rect 10961 7110 13327 7112
rect 10961 7107 11027 7110
rect 12801 7107 12867 7110
rect 13261 7107 13327 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 5993 7034 6059 7037
rect 6361 7034 6427 7037
rect 8334 7034 8340 7036
rect 5993 7032 8340 7034
rect 5993 6976 5998 7032
rect 6054 6976 6366 7032
rect 6422 6976 8340 7032
rect 5993 6974 8340 6976
rect 5993 6971 6059 6974
rect 6361 6971 6427 6974
rect 8334 6972 8340 6974
rect 8404 6972 8410 7036
rect 7925 6900 7991 6901
rect 7925 6896 7972 6900
rect 8036 6898 8042 6900
rect 7925 6840 7930 6896
rect 7925 6836 7972 6840
rect 8036 6838 8082 6898
rect 12065 6896 12131 6901
rect 15285 6900 15351 6901
rect 15285 6898 15332 6900
rect 12065 6840 12070 6896
rect 12126 6840 12131 6896
rect 8036 6836 8042 6838
rect 7925 6835 7991 6836
rect 12065 6835 12131 6840
rect 15240 6896 15332 6898
rect 15240 6840 15290 6896
rect 15240 6838 15332 6840
rect 15285 6836 15332 6838
rect 15396 6836 15402 6900
rect 15285 6835 15351 6836
rect 5717 6764 5783 6765
rect 5717 6762 5764 6764
rect 5672 6760 5764 6762
rect 5672 6704 5722 6760
rect 5672 6702 5764 6704
rect 5717 6700 5764 6702
rect 5828 6700 5834 6764
rect 11789 6762 11855 6765
rect 12068 6762 12128 6835
rect 11789 6760 12128 6762
rect 11789 6704 11794 6760
rect 11850 6704 12128 6760
rect 11789 6702 12128 6704
rect 5717 6699 5783 6700
rect 11789 6699 11855 6702
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 7557 6490 7623 6493
rect 7833 6490 7899 6493
rect 7557 6488 7899 6490
rect 7557 6432 7562 6488
rect 7618 6432 7838 6488
rect 7894 6432 7899 6488
rect 7557 6430 7899 6432
rect 7557 6427 7623 6430
rect 7833 6427 7899 6430
rect 10777 6490 10843 6493
rect 13353 6490 13419 6493
rect 10777 6488 13419 6490
rect 10777 6432 10782 6488
rect 10838 6432 13358 6488
rect 13414 6432 13419 6488
rect 10777 6430 13419 6432
rect 10777 6427 10843 6430
rect 13353 6427 13419 6430
rect 3366 6292 3372 6356
rect 3436 6354 3442 6356
rect 3509 6354 3575 6357
rect 3436 6352 3575 6354
rect 3436 6296 3514 6352
rect 3570 6296 3575 6352
rect 3436 6294 3575 6296
rect 3436 6292 3442 6294
rect 3509 6291 3575 6294
rect 3693 6354 3759 6357
rect 4889 6354 4955 6357
rect 6453 6354 6519 6357
rect 3693 6352 6519 6354
rect 3693 6296 3698 6352
rect 3754 6296 4894 6352
rect 4950 6296 6458 6352
rect 6514 6296 6519 6352
rect 3693 6294 6519 6296
rect 3693 6291 3759 6294
rect 4889 6291 4955 6294
rect 6453 6291 6519 6294
rect 10409 6354 10475 6357
rect 11329 6354 11395 6357
rect 10409 6352 11395 6354
rect 10409 6296 10414 6352
rect 10470 6296 11334 6352
rect 11390 6296 11395 6352
rect 10409 6294 11395 6296
rect 10409 6291 10475 6294
rect 11329 6291 11395 6294
rect 13302 6292 13308 6356
rect 13372 6354 13378 6356
rect 14273 6354 14339 6357
rect 13372 6352 14339 6354
rect 13372 6296 14278 6352
rect 14334 6296 14339 6352
rect 13372 6294 14339 6296
rect 13372 6292 13378 6294
rect 14273 6291 14339 6294
rect 3182 6156 3188 6220
rect 3252 6218 3258 6220
rect 4797 6218 4863 6221
rect 3252 6216 4863 6218
rect 3252 6160 4802 6216
rect 4858 6160 4863 6216
rect 3252 6158 4863 6160
rect 3252 6156 3258 6158
rect 4797 6155 4863 6158
rect 8753 6218 8819 6221
rect 9581 6218 9647 6221
rect 8753 6216 9647 6218
rect 8753 6160 8758 6216
rect 8814 6160 9586 6216
rect 9642 6160 9647 6216
rect 8753 6158 9647 6160
rect 8753 6155 8819 6158
rect 9581 6155 9647 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 7373 5946 7439 5949
rect 4662 5944 7439 5946
rect 4662 5888 7378 5944
rect 7434 5888 7439 5944
rect 4662 5886 7439 5888
rect 3601 5810 3667 5813
rect 4662 5810 4722 5886
rect 7373 5883 7439 5886
rect 7741 5946 7807 5949
rect 12157 5946 12223 5949
rect 14917 5946 14983 5949
rect 7741 5944 14983 5946
rect 7741 5888 7746 5944
rect 7802 5888 12162 5944
rect 12218 5888 14922 5944
rect 14978 5888 14983 5944
rect 7741 5886 14983 5888
rect 7741 5883 7807 5886
rect 12157 5883 12223 5886
rect 14917 5883 14983 5886
rect 3601 5808 4722 5810
rect 3601 5752 3606 5808
rect 3662 5752 4722 5808
rect 3601 5750 4722 5752
rect 8477 5810 8543 5813
rect 10317 5810 10383 5813
rect 12065 5810 12131 5813
rect 13629 5812 13695 5813
rect 13629 5810 13676 5812
rect 8477 5808 12131 5810
rect 8477 5752 8482 5808
rect 8538 5752 10322 5808
rect 10378 5752 12070 5808
rect 12126 5752 12131 5808
rect 8477 5750 12131 5752
rect 13584 5808 13676 5810
rect 13584 5752 13634 5808
rect 13584 5750 13676 5752
rect 3601 5747 3667 5750
rect 8477 5747 8543 5750
rect 10317 5747 10383 5750
rect 12065 5747 12131 5750
rect 13629 5748 13676 5750
rect 13740 5748 13746 5812
rect 13629 5747 13695 5748
rect 3049 5674 3115 5677
rect 12985 5674 13051 5677
rect 3049 5672 13051 5674
rect 3049 5616 3054 5672
rect 3110 5616 12990 5672
rect 13046 5616 13051 5672
rect 3049 5614 13051 5616
rect 3049 5611 3115 5614
rect 12985 5611 13051 5614
rect 14222 5612 14228 5676
rect 14292 5674 14298 5676
rect 14365 5674 14431 5677
rect 14292 5672 14431 5674
rect 14292 5616 14370 5672
rect 14426 5616 14431 5672
rect 14292 5614 14431 5616
rect 14292 5612 14298 5614
rect 14365 5611 14431 5614
rect 0 5538 800 5568
rect 1485 5538 1551 5541
rect 0 5536 1551 5538
rect 0 5480 1490 5536
rect 1546 5480 1551 5536
rect 0 5478 1551 5480
rect 0 5448 800 5478
rect 1485 5475 1551 5478
rect 6913 5538 6979 5541
rect 7414 5538 7420 5540
rect 6913 5536 7420 5538
rect 6913 5480 6918 5536
rect 6974 5480 7420 5536
rect 6913 5478 7420 5480
rect 6913 5475 6979 5478
rect 7414 5476 7420 5478
rect 7484 5476 7490 5540
rect 10593 5538 10659 5541
rect 14273 5538 14339 5541
rect 10593 5536 14339 5538
rect 10593 5480 10598 5536
rect 10654 5480 14278 5536
rect 14334 5480 14339 5536
rect 10593 5478 14339 5480
rect 10593 5475 10659 5478
rect 14273 5475 14339 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 5901 5402 5967 5405
rect 8845 5402 8911 5405
rect 9489 5402 9555 5405
rect 5901 5400 9555 5402
rect 5901 5344 5906 5400
rect 5962 5344 8850 5400
rect 8906 5344 9494 5400
rect 9550 5344 9555 5400
rect 5901 5342 9555 5344
rect 5901 5339 5967 5342
rect 8845 5339 8911 5342
rect 9489 5339 9555 5342
rect 8845 5268 8911 5269
rect 8845 5266 8892 5268
rect 8800 5264 8892 5266
rect 8800 5208 8850 5264
rect 8800 5206 8892 5208
rect 8845 5204 8892 5206
rect 8956 5204 8962 5268
rect 8845 5203 8911 5204
rect 11973 4994 12039 4997
rect 13629 4994 13695 4997
rect 11973 4992 13695 4994
rect 11973 4936 11978 4992
rect 12034 4936 13634 4992
rect 13690 4936 13695 4992
rect 11973 4934 13695 4936
rect 11973 4931 12039 4934
rect 13629 4931 13695 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 5349 4586 5415 4589
rect 12014 4586 12020 4588
rect 5349 4584 12020 4586
rect 5349 4528 5354 4584
rect 5410 4528 12020 4584
rect 5349 4526 12020 4528
rect 5349 4523 5415 4526
rect 12014 4524 12020 4526
rect 12084 4586 12090 4588
rect 13169 4586 13235 4589
rect 12084 4584 13235 4586
rect 12084 4528 13174 4584
rect 13230 4528 13235 4584
rect 12084 4526 13235 4528
rect 12084 4524 12090 4526
rect 13169 4523 13235 4526
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 10593 4178 10659 4181
rect 14774 4178 14780 4180
rect 10593 4176 14780 4178
rect 10593 4120 10598 4176
rect 10654 4120 14780 4176
rect 10593 4118 14780 4120
rect 10593 4115 10659 4118
rect 14774 4116 14780 4118
rect 14844 4116 14850 4180
rect 6862 3980 6868 4044
rect 6932 4042 6938 4044
rect 7005 4042 7071 4045
rect 6932 4040 7071 4042
rect 6932 3984 7010 4040
rect 7066 3984 7071 4040
rect 6932 3982 7071 3984
rect 6932 3980 6938 3982
rect 7005 3979 7071 3982
rect 13261 4042 13327 4045
rect 13486 4042 13492 4044
rect 13261 4040 13492 4042
rect 13261 3984 13266 4040
rect 13322 3984 13492 4040
rect 13261 3982 13492 3984
rect 13261 3979 13327 3982
rect 13486 3980 13492 3982
rect 13556 3980 13562 4044
rect 9581 3906 9647 3909
rect 13302 3906 13308 3908
rect 9581 3904 13308 3906
rect 9581 3848 9586 3904
rect 9642 3848 13308 3904
rect 9581 3846 13308 3848
rect 9581 3843 9647 3846
rect 13302 3844 13308 3846
rect 13372 3906 13378 3908
rect 13721 3906 13787 3909
rect 13372 3904 13787 3906
rect 13372 3848 13726 3904
rect 13782 3848 13787 3904
rect 13372 3846 13787 3848
rect 13372 3844 13378 3846
rect 13721 3843 13787 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 12198 3572 12204 3636
rect 12268 3634 12274 3636
rect 13077 3634 13143 3637
rect 12268 3632 13143 3634
rect 12268 3576 13082 3632
rect 13138 3576 13143 3632
rect 12268 3574 13143 3576
rect 12268 3572 12274 3574
rect 13077 3571 13143 3574
rect 2773 3498 2839 3501
rect 9949 3498 10015 3501
rect 10174 3498 10180 3500
rect 2773 3496 10180 3498
rect 2773 3440 2778 3496
rect 2834 3440 9954 3496
rect 10010 3440 10180 3496
rect 2773 3438 10180 3440
rect 2773 3435 2839 3438
rect 9949 3435 10015 3438
rect 10174 3436 10180 3438
rect 10244 3498 10250 3500
rect 10685 3498 10751 3501
rect 10244 3496 10751 3498
rect 10244 3440 10690 3496
rect 10746 3440 10751 3496
rect 10244 3438 10751 3440
rect 10244 3436 10250 3438
rect 10685 3435 10751 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 8661 3090 8727 3093
rect 12709 3090 12775 3093
rect 8661 3088 12775 3090
rect 8661 3032 8666 3088
rect 8722 3032 12714 3088
rect 12770 3032 12775 3088
rect 8661 3030 12775 3032
rect 8661 3027 8727 3030
rect 12709 3027 12775 3030
rect 6361 2954 6427 2957
rect 10317 2954 10383 2957
rect 6361 2952 10383 2954
rect 6361 2896 6366 2952
rect 6422 2896 10322 2952
rect 10378 2896 10383 2952
rect 6361 2894 10383 2896
rect 6361 2891 6427 2894
rect 10317 2891 10383 2894
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 5580 16492 5644 16556
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 9260 16008 9324 16012
rect 9260 15952 9310 16008
rect 9310 15952 9324 16008
rect 9260 15948 9324 15952
rect 8892 15872 8956 15876
rect 8892 15816 8942 15872
rect 8942 15816 8956 15872
rect 8892 15812 8956 15816
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 6684 15676 6748 15740
rect 4660 15464 4724 15468
rect 4660 15408 4674 15464
rect 4674 15408 4724 15464
rect 4660 15404 4724 15408
rect 14780 15404 14844 15468
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 9628 14996 9692 15060
rect 9444 14920 9508 14924
rect 9444 14864 9458 14920
rect 9458 14864 9508 14920
rect 9444 14860 9508 14864
rect 7972 14724 8036 14788
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 15516 14452 15580 14516
rect 3924 14316 3988 14380
rect 12388 14316 12452 14380
rect 7052 14180 7116 14244
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 6132 14044 6196 14108
rect 4660 13908 4724 13972
rect 6500 13772 6564 13836
rect 9812 13772 9876 13836
rect 16068 13832 16132 13836
rect 16068 13776 16082 13832
rect 16082 13776 16132 13832
rect 16068 13772 16132 13776
rect 16436 13772 16500 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 3188 13288 3252 13292
rect 3188 13232 3202 13288
rect 3202 13232 3252 13288
rect 3188 13228 3252 13232
rect 12572 13228 12636 13292
rect 11284 13152 11348 13156
rect 11284 13096 11334 13152
rect 11334 13096 11348 13152
rect 11284 13092 11348 13096
rect 11652 13092 11716 13156
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 5764 12684 5828 12748
rect 3004 12608 3068 12612
rect 3004 12552 3054 12608
rect 3054 12552 3068 12608
rect 3004 12548 3068 12552
rect 7420 12684 7484 12748
rect 15148 12684 15212 12748
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 7236 12412 7300 12476
rect 9076 12412 9140 12476
rect 5396 12140 5460 12204
rect 14412 12200 14476 12204
rect 14412 12144 14426 12200
rect 14426 12144 14476 12200
rect 14412 12140 14476 12144
rect 14964 12200 15028 12204
rect 14964 12144 15014 12200
rect 15014 12144 15028 12200
rect 14964 12140 15028 12144
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 8340 11868 8404 11932
rect 15332 11732 15396 11796
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 6868 11248 6932 11252
rect 6868 11192 6918 11248
rect 6918 11192 6932 11248
rect 6868 11188 6932 11192
rect 11284 11188 11348 11252
rect 6684 11052 6748 11116
rect 10916 11052 10980 11116
rect 13308 11052 13372 11116
rect 8340 10916 8404 10980
rect 11652 10916 11716 10980
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 6500 10780 6564 10844
rect 13492 10644 13556 10708
rect 14964 10704 15028 10708
rect 14964 10648 14978 10704
rect 14978 10648 15028 10704
rect 14964 10644 15028 10648
rect 15148 10644 15212 10708
rect 4660 10508 4724 10572
rect 12388 10508 12452 10572
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 9076 10236 9140 10300
rect 3924 9964 3988 10028
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 3372 9752 3436 9756
rect 3372 9696 3386 9752
rect 3386 9696 3436 9752
rect 3372 9692 3436 9696
rect 12020 9692 12084 9756
rect 3004 9616 3068 9620
rect 3004 9560 3054 9616
rect 3054 9560 3068 9616
rect 3004 9556 3068 9560
rect 6132 9556 6196 9620
rect 7236 9556 7300 9620
rect 14412 9556 14476 9620
rect 16436 9616 16500 9620
rect 16436 9560 16486 9616
rect 16486 9560 16500 9616
rect 16436 9556 16500 9560
rect 5580 9420 5644 9484
rect 9628 9420 9692 9484
rect 14228 9420 14292 9484
rect 16068 9344 16132 9348
rect 16068 9288 16118 9344
rect 16118 9288 16132 9344
rect 16068 9284 16132 9288
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 7052 9012 7116 9076
rect 3004 8876 3068 8940
rect 6684 8876 6748 8940
rect 14780 8876 14844 8940
rect 7236 8740 7300 8804
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 15516 8468 15580 8532
rect 9260 8196 9324 8260
rect 9812 8196 9876 8260
rect 13676 8332 13740 8396
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 9444 7924 9508 7988
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 10916 7380 10980 7444
rect 5396 7304 5460 7308
rect 5396 7248 5410 7304
rect 5410 7248 5460 7304
rect 5396 7244 5460 7248
rect 10180 7244 10244 7308
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 8340 6972 8404 7036
rect 7972 6896 8036 6900
rect 7972 6840 7986 6896
rect 7986 6840 8036 6896
rect 7972 6836 8036 6840
rect 15332 6896 15396 6900
rect 15332 6840 15346 6896
rect 15346 6840 15396 6896
rect 15332 6836 15396 6840
rect 5764 6760 5828 6764
rect 5764 6704 5778 6760
rect 5778 6704 5828 6760
rect 5764 6700 5828 6704
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 3372 6292 3436 6356
rect 13308 6292 13372 6356
rect 3188 6156 3252 6220
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 13676 5808 13740 5812
rect 13676 5752 13690 5808
rect 13690 5752 13740 5808
rect 13676 5748 13740 5752
rect 14228 5612 14292 5676
rect 7420 5476 7484 5540
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 8892 5264 8956 5268
rect 8892 5208 8906 5264
rect 8906 5208 8956 5264
rect 8892 5204 8956 5208
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 12020 4524 12084 4588
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 14780 4116 14844 4180
rect 6868 3980 6932 4044
rect 13492 3980 13556 4044
rect 13308 3844 13372 3908
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 12204 3572 12268 3636
rect 10180 3436 10244 3500
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 19072 4528 19088
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4868 18528 5188 19088
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 5579 16556 5645 16557
rect 5579 16492 5580 16556
rect 5644 16492 5645 16556
rect 5579 16491 5645 16492
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4659 15468 4725 15469
rect 4659 15404 4660 15468
rect 4724 15404 4725 15468
rect 4659 15403 4725 15404
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 3923 14380 3989 14381
rect 3923 14316 3924 14380
rect 3988 14316 3989 14380
rect 3923 14315 3989 14316
rect 3187 13292 3253 13293
rect 3187 13228 3188 13292
rect 3252 13228 3253 13292
rect 3187 13227 3253 13228
rect 3003 12612 3069 12613
rect 3003 12548 3004 12612
rect 3068 12548 3069 12612
rect 3003 12547 3069 12548
rect 3006 9621 3066 12547
rect 3003 9620 3069 9621
rect 3003 9556 3004 9620
rect 3068 9556 3069 9620
rect 3003 9555 3069 9556
rect 3006 8941 3066 9555
rect 3003 8940 3069 8941
rect 3003 8876 3004 8940
rect 3068 8876 3069 8940
rect 3003 8875 3069 8876
rect 3190 6221 3250 13227
rect 3926 10029 3986 14315
rect 4208 13632 4528 14656
rect 4662 13973 4722 15403
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4659 13972 4725 13973
rect 4659 13908 4660 13972
rect 4724 13908 4725 13972
rect 4659 13907 4725 13908
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4662 10573 4722 13907
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 5395 12204 5461 12205
rect 5395 12140 5396 12204
rect 5460 12140 5461 12204
rect 5395 12139 5461 12140
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4659 10572 4725 10573
rect 4659 10508 4660 10572
rect 4724 10508 4725 10572
rect 4659 10507 4725 10508
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 3923 10028 3989 10029
rect 3923 9964 3924 10028
rect 3988 9964 3989 10028
rect 3923 9963 3989 9964
rect 3371 9756 3437 9757
rect 3371 9692 3372 9756
rect 3436 9692 3437 9756
rect 3371 9691 3437 9692
rect 3374 6357 3434 9691
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 3371 6356 3437 6357
rect 3371 6292 3372 6356
rect 3436 6292 3437 6356
rect 3371 6291 3437 6292
rect 3187 6220 3253 6221
rect 3187 6156 3188 6220
rect 3252 6156 3253 6220
rect 3187 6155 3253 6156
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 5398 7309 5458 12139
rect 5582 9485 5642 16491
rect 9259 16012 9325 16013
rect 9259 15948 9260 16012
rect 9324 15948 9325 16012
rect 9259 15947 9325 15948
rect 8891 15876 8957 15877
rect 8891 15812 8892 15876
rect 8956 15812 8957 15876
rect 8891 15811 8957 15812
rect 6683 15740 6749 15741
rect 6683 15676 6684 15740
rect 6748 15676 6749 15740
rect 6683 15675 6749 15676
rect 6131 14108 6197 14109
rect 6131 14044 6132 14108
rect 6196 14044 6197 14108
rect 6131 14043 6197 14044
rect 5763 12748 5829 12749
rect 5763 12684 5764 12748
rect 5828 12684 5829 12748
rect 5763 12683 5829 12684
rect 5579 9484 5645 9485
rect 5579 9420 5580 9484
rect 5644 9420 5645 9484
rect 5579 9419 5645 9420
rect 5395 7308 5461 7309
rect 5395 7244 5396 7308
rect 5460 7244 5461 7308
rect 5395 7243 5461 7244
rect 5766 6765 5826 12683
rect 6134 9621 6194 14043
rect 6499 13836 6565 13837
rect 6499 13772 6500 13836
rect 6564 13772 6565 13836
rect 6499 13771 6565 13772
rect 6502 10845 6562 13771
rect 6686 11117 6746 15675
rect 7971 14788 8037 14789
rect 7971 14724 7972 14788
rect 8036 14724 8037 14788
rect 7971 14723 8037 14724
rect 7051 14244 7117 14245
rect 7051 14180 7052 14244
rect 7116 14180 7117 14244
rect 7051 14179 7117 14180
rect 6867 11252 6933 11253
rect 6867 11188 6868 11252
rect 6932 11188 6933 11252
rect 6867 11187 6933 11188
rect 6683 11116 6749 11117
rect 6683 11052 6684 11116
rect 6748 11052 6749 11116
rect 6683 11051 6749 11052
rect 6499 10844 6565 10845
rect 6499 10780 6500 10844
rect 6564 10780 6565 10844
rect 6499 10779 6565 10780
rect 6131 9620 6197 9621
rect 6131 9556 6132 9620
rect 6196 9556 6197 9620
rect 6131 9555 6197 9556
rect 6686 8941 6746 11051
rect 6683 8940 6749 8941
rect 6683 8876 6684 8940
rect 6748 8876 6749 8940
rect 6683 8875 6749 8876
rect 5763 6764 5829 6765
rect 5763 6700 5764 6764
rect 5828 6700 5829 6764
rect 5763 6699 5829 6700
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 6870 4045 6930 11187
rect 7054 9077 7114 14179
rect 7419 12748 7485 12749
rect 7419 12684 7420 12748
rect 7484 12684 7485 12748
rect 7419 12683 7485 12684
rect 7235 12476 7301 12477
rect 7235 12412 7236 12476
rect 7300 12412 7301 12476
rect 7235 12411 7301 12412
rect 7238 9621 7298 12411
rect 7235 9620 7301 9621
rect 7235 9556 7236 9620
rect 7300 9556 7301 9620
rect 7235 9555 7301 9556
rect 7051 9076 7117 9077
rect 7051 9012 7052 9076
rect 7116 9012 7117 9076
rect 7051 9011 7117 9012
rect 7238 8805 7298 9555
rect 7235 8804 7301 8805
rect 7235 8740 7236 8804
rect 7300 8740 7301 8804
rect 7235 8739 7301 8740
rect 7422 5541 7482 12683
rect 7974 6901 8034 14723
rect 8339 11932 8405 11933
rect 8339 11868 8340 11932
rect 8404 11868 8405 11932
rect 8339 11867 8405 11868
rect 8342 10981 8402 11867
rect 8339 10980 8405 10981
rect 8339 10916 8340 10980
rect 8404 10916 8405 10980
rect 8339 10915 8405 10916
rect 8342 7037 8402 10915
rect 8339 7036 8405 7037
rect 8339 6972 8340 7036
rect 8404 6972 8405 7036
rect 8339 6971 8405 6972
rect 7971 6900 8037 6901
rect 7971 6836 7972 6900
rect 8036 6836 8037 6900
rect 7971 6835 8037 6836
rect 7419 5540 7485 5541
rect 7419 5476 7420 5540
rect 7484 5476 7485 5540
rect 7419 5475 7485 5476
rect 8894 5269 8954 15811
rect 9075 12476 9141 12477
rect 9075 12412 9076 12476
rect 9140 12412 9141 12476
rect 9075 12411 9141 12412
rect 9078 10301 9138 12411
rect 9075 10300 9141 10301
rect 9075 10236 9076 10300
rect 9140 10236 9141 10300
rect 9075 10235 9141 10236
rect 9262 8261 9322 15947
rect 14779 15468 14845 15469
rect 14779 15404 14780 15468
rect 14844 15404 14845 15468
rect 14779 15403 14845 15404
rect 9627 15060 9693 15061
rect 9627 14996 9628 15060
rect 9692 14996 9693 15060
rect 9627 14995 9693 14996
rect 9443 14924 9509 14925
rect 9443 14860 9444 14924
rect 9508 14860 9509 14924
rect 9443 14859 9509 14860
rect 9259 8260 9325 8261
rect 9259 8196 9260 8260
rect 9324 8196 9325 8260
rect 9259 8195 9325 8196
rect 9446 7989 9506 14859
rect 9630 9485 9690 14995
rect 12387 14380 12453 14381
rect 12387 14316 12388 14380
rect 12452 14316 12453 14380
rect 12387 14315 12453 14316
rect 9811 13836 9877 13837
rect 9811 13772 9812 13836
rect 9876 13772 9877 13836
rect 9811 13771 9877 13772
rect 9627 9484 9693 9485
rect 9627 9420 9628 9484
rect 9692 9420 9693 9484
rect 9627 9419 9693 9420
rect 9814 8261 9874 13771
rect 11283 13156 11349 13157
rect 11283 13092 11284 13156
rect 11348 13092 11349 13156
rect 11283 13091 11349 13092
rect 11651 13156 11717 13157
rect 11651 13092 11652 13156
rect 11716 13092 11717 13156
rect 11651 13091 11717 13092
rect 11286 11253 11346 13091
rect 11283 11252 11349 11253
rect 11283 11188 11284 11252
rect 11348 11188 11349 11252
rect 11283 11187 11349 11188
rect 10915 11116 10981 11117
rect 10915 11052 10916 11116
rect 10980 11052 10981 11116
rect 10915 11051 10981 11052
rect 9811 8260 9877 8261
rect 9811 8196 9812 8260
rect 9876 8196 9877 8260
rect 9811 8195 9877 8196
rect 9443 7988 9509 7989
rect 9443 7924 9444 7988
rect 9508 7924 9509 7988
rect 9443 7923 9509 7924
rect 10918 7445 10978 11051
rect 11654 10981 11714 13091
rect 11651 10980 11717 10981
rect 11651 10916 11652 10980
rect 11716 10916 11717 10980
rect 11651 10915 11717 10916
rect 12390 10573 12450 14315
rect 12571 13292 12637 13293
rect 12571 13228 12572 13292
rect 12636 13228 12637 13292
rect 12571 13227 12637 13228
rect 12387 10572 12453 10573
rect 12387 10508 12388 10572
rect 12452 10508 12453 10572
rect 12387 10507 12453 10508
rect 12019 9756 12085 9757
rect 12019 9692 12020 9756
rect 12084 9692 12085 9756
rect 12019 9691 12085 9692
rect 10915 7444 10981 7445
rect 10915 7380 10916 7444
rect 10980 7380 10981 7444
rect 10915 7379 10981 7380
rect 10179 7308 10245 7309
rect 10179 7244 10180 7308
rect 10244 7244 10245 7308
rect 10179 7243 10245 7244
rect 8891 5268 8957 5269
rect 8891 5204 8892 5268
rect 8956 5204 8957 5268
rect 8891 5203 8957 5204
rect 6867 4044 6933 4045
rect 6867 3980 6868 4044
rect 6932 3980 6933 4044
rect 6867 3979 6933 3980
rect 10182 3501 10242 7243
rect 12022 4589 12082 9691
rect 12574 6930 12634 13227
rect 14411 12204 14477 12205
rect 14411 12140 14412 12204
rect 14476 12140 14477 12204
rect 14411 12139 14477 12140
rect 13307 11116 13373 11117
rect 13307 11052 13308 11116
rect 13372 11052 13373 11116
rect 13307 11051 13373 11052
rect 12206 6870 12634 6930
rect 12019 4588 12085 4589
rect 12019 4524 12020 4588
rect 12084 4524 12085 4588
rect 12019 4523 12085 4524
rect 12206 3637 12266 6870
rect 13310 6357 13370 11051
rect 13491 10708 13557 10709
rect 13491 10644 13492 10708
rect 13556 10644 13557 10708
rect 13491 10643 13557 10644
rect 13307 6356 13373 6357
rect 13307 6292 13308 6356
rect 13372 6292 13373 6356
rect 13307 6291 13373 6292
rect 13310 3909 13370 6291
rect 13494 4045 13554 10643
rect 14414 9621 14474 12139
rect 14411 9620 14477 9621
rect 14411 9556 14412 9620
rect 14476 9556 14477 9620
rect 14411 9555 14477 9556
rect 14227 9484 14293 9485
rect 14227 9420 14228 9484
rect 14292 9420 14293 9484
rect 14227 9419 14293 9420
rect 13675 8396 13741 8397
rect 13675 8332 13676 8396
rect 13740 8332 13741 8396
rect 13675 8331 13741 8332
rect 13678 5813 13738 8331
rect 13675 5812 13741 5813
rect 13675 5748 13676 5812
rect 13740 5748 13741 5812
rect 13675 5747 13741 5748
rect 14230 5677 14290 9419
rect 14782 8941 14842 15403
rect 15515 14516 15581 14517
rect 15515 14452 15516 14516
rect 15580 14452 15581 14516
rect 15515 14451 15581 14452
rect 15147 12748 15213 12749
rect 15147 12684 15148 12748
rect 15212 12684 15213 12748
rect 15147 12683 15213 12684
rect 14963 12204 15029 12205
rect 14963 12140 14964 12204
rect 15028 12140 15029 12204
rect 14963 12139 15029 12140
rect 14966 10709 15026 12139
rect 15150 10709 15210 12683
rect 15331 11796 15397 11797
rect 15331 11732 15332 11796
rect 15396 11732 15397 11796
rect 15331 11731 15397 11732
rect 14963 10708 15029 10709
rect 14963 10644 14964 10708
rect 15028 10644 15029 10708
rect 14963 10643 15029 10644
rect 15147 10708 15213 10709
rect 15147 10644 15148 10708
rect 15212 10644 15213 10708
rect 15147 10643 15213 10644
rect 14779 8940 14845 8941
rect 14779 8876 14780 8940
rect 14844 8876 14845 8940
rect 14779 8875 14845 8876
rect 14227 5676 14293 5677
rect 14227 5612 14228 5676
rect 14292 5612 14293 5676
rect 14227 5611 14293 5612
rect 14782 4181 14842 8875
rect 15334 6901 15394 11731
rect 15518 8533 15578 14451
rect 16067 13836 16133 13837
rect 16067 13772 16068 13836
rect 16132 13772 16133 13836
rect 16067 13771 16133 13772
rect 16435 13836 16501 13837
rect 16435 13772 16436 13836
rect 16500 13772 16501 13836
rect 16435 13771 16501 13772
rect 16070 9349 16130 13771
rect 16438 9621 16498 13771
rect 16435 9620 16501 9621
rect 16435 9556 16436 9620
rect 16500 9556 16501 9620
rect 16435 9555 16501 9556
rect 16067 9348 16133 9349
rect 16067 9284 16068 9348
rect 16132 9284 16133 9348
rect 16067 9283 16133 9284
rect 15515 8532 15581 8533
rect 15515 8468 15516 8532
rect 15580 8468 15581 8532
rect 15515 8467 15581 8468
rect 15331 6900 15397 6901
rect 15331 6836 15332 6900
rect 15396 6836 15397 6900
rect 15331 6835 15397 6836
rect 14779 4180 14845 4181
rect 14779 4116 14780 4180
rect 14844 4116 14845 4180
rect 14779 4115 14845 4116
rect 13491 4044 13557 4045
rect 13491 3980 13492 4044
rect 13556 3980 13557 4044
rect 13491 3979 13557 3980
rect 13307 3908 13373 3909
rect 13307 3844 13308 3908
rect 13372 3844 13373 3908
rect 13307 3843 13373 3844
rect 12203 3636 12269 3637
rect 12203 3572 12204 3636
rect 12268 3572 12269 3636
rect 12203 3571 12269 3572
rect 10179 3500 10245 3501
rect 10179 3436 10180 3500
rect 10244 3436 10245 3500
rect 10179 3435 10245 3436
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _391_
timestamp 1
transform -1 0 16376 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp 1
transform 1 0 10580 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 1
transform 1 0 5888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp 1
transform -1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _395_
timestamp 1
transform -1 0 16560 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _396_
timestamp 1
transform 1 0 7728 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _397_
timestamp 1
transform 1 0 2576 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp 1
transform -1 0 17388 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _399_
timestamp 1
transform 1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _400_
timestamp 1
transform 1 0 7912 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _401_
timestamp 1
transform -1 0 17112 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _402_
timestamp 1
transform -1 0 2852 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _403_
timestamp 1
transform 1 0 16652 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp 1
transform 1 0 15916 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _405_
timestamp 1
transform -1 0 5888 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _406_
timestamp 1
transform -1 0 11040 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _407_
timestamp 1
transform 1 0 4048 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _408_
timestamp 1
transform 1 0 6440 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _409_
timestamp 1
transform 1 0 2944 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _410_
timestamp 1
transform -1 0 13616 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _411_
timestamp 1
transform 1 0 4692 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _412_
timestamp 1
transform 1 0 2300 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _413_
timestamp 1
transform -1 0 6992 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _414_
timestamp 1
transform 1 0 1932 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _415_
timestamp 1
transform -1 0 14536 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _416_
timestamp 1
transform -1 0 14812 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _417_
timestamp 1
transform 1 0 3220 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _418_
timestamp 1
transform 1 0 2668 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__o21ai_4  _419_
timestamp 1
transform 1 0 5520 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _420_
timestamp 1
transform -1 0 8740 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _421_
timestamp 1
transform 1 0 3772 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _422_
timestamp 1
transform 1 0 5980 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_1  _423_
timestamp 1
transform 1 0 11868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _424_
timestamp 1
transform 1 0 11868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _425_
timestamp 1
transform -1 0 15732 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _426_
timestamp 1
transform -1 0 16560 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _427_
timestamp 1
transform 1 0 14996 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _428_
timestamp 1
transform -1 0 13340 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _429_
timestamp 1
transform 1 0 6348 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_4  _430_
timestamp 1
transform -1 0 16744 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__and2_1  _431_
timestamp 1
transform -1 0 10396 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _432_
timestamp 1
transform -1 0 10304 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _433_
timestamp 1
transform 1 0 8924 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _434_
timestamp 1
transform 1 0 4968 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _435_
timestamp 1
transform -1 0 12328 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _436_
timestamp 1
transform -1 0 11316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _437_
timestamp 1
transform 1 0 10672 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_2  _438_
timestamp 1
transform 1 0 16560 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _439_
timestamp 1
transform -1 0 13524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _440_
timestamp 1
transform 1 0 11316 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _441_
timestamp 1
transform -1 0 11868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _442_
timestamp 1
transform 1 0 2852 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _443_
timestamp 1
transform -1 0 5428 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _444_
timestamp 1
transform -1 0 8832 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _445_
timestamp 1
transform -1 0 9200 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _446_
timestamp 1
transform -1 0 12328 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _447_
timestamp 1
transform -1 0 12512 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _448_
timestamp 1
transform -1 0 17848 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _449_
timestamp 1
transform 1 0 10396 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _450_
timestamp 1
transform 1 0 9660 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_2  _451_
timestamp 1
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_2  _452_
timestamp 1
transform -1 0 8004 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _453_
timestamp 1
transform 1 0 9108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _454_
timestamp 1
transform -1 0 16928 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _455_
timestamp 1
transform -1 0 5428 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _456_
timestamp 1
transform 1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _457_
timestamp 1
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _458_
timestamp 1
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _459_
timestamp 1
transform 1 0 2668 0 -1 4352
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _460_
timestamp 1
transform 1 0 9936 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _461_
timestamp 1
transform 1 0 11684 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _462_
timestamp 1
transform 1 0 5244 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _463_
timestamp 1
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _464_
timestamp 1
transform -1 0 7176 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _465_
timestamp 1
transform 1 0 14996 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _466_
timestamp 1
transform -1 0 9752 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _467_
timestamp 1
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _468_
timestamp 1
transform 1 0 9844 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _469_
timestamp 1
transform -1 0 16376 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_2  _470_
timestamp 1
transform 1 0 16652 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _471_
timestamp 1
transform 1 0 17296 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _472_
timestamp 1
transform -1 0 9660 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _473_
timestamp 1
transform -1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _474_
timestamp 1
transform -1 0 9016 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _475_
timestamp 1
transform 1 0 4968 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _476_
timestamp 1
transform -1 0 15732 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _477_
timestamp 1
transform -1 0 8648 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _478_
timestamp 1
transform 1 0 5520 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_4  _479_
timestamp 1
transform 1 0 2208 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__nor2_1  _480_
timestamp 1
transform 1 0 2944 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _481_
timestamp 1
transform 1 0 2760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _482_
timestamp 1
transform 1 0 3772 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _483_
timestamp 1
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _484_
timestamp 1
transform -1 0 7728 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _485_
timestamp 1
transform 1 0 10488 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _486_
timestamp 1
transform -1 0 8096 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _487_
timestamp 1
transform -1 0 7636 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _488_
timestamp 1
transform -1 0 8556 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _489_
timestamp 1
transform 1 0 9292 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _490_
timestamp 1
transform 1 0 10028 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _491_
timestamp 1
transform -1 0 16560 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _492_
timestamp 1
transform -1 0 10212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _493_
timestamp 1
transform -1 0 5152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _494_
timestamp 1
transform -1 0 4968 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _495_
timestamp 1
transform -1 0 12972 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_1  _496_
timestamp 1
transform 1 0 9752 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _497_
timestamp 1
transform -1 0 10396 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _498_
timestamp 1
transform -1 0 14444 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _499_
timestamp 1
transform 1 0 11776 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _500_
timestamp 1
transform 1 0 14812 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _501_
timestamp 1
transform 1 0 6992 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _502_
timestamp 1
transform 1 0 12236 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _503_
timestamp 1
transform -1 0 5888 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _504_
timestamp 1
transform 1 0 3312 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _505_
timestamp 1
transform -1 0 4324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _506_
timestamp 1
transform 1 0 4416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _507_
timestamp 1
transform 1 0 5336 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _508_
timestamp 1
transform 1 0 5060 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _509_
timestamp 1
transform -1 0 6348 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _510_
timestamp 1
transform -1 0 7360 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_4  _511_
timestamp 1
transform 1 0 14812 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _512_
timestamp 1
transform -1 0 7636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _513_
timestamp 1
transform 1 0 6992 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _514_
timestamp 1
transform 1 0 5796 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _515_
timestamp 1
transform -1 0 8004 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _516_
timestamp 1
transform 1 0 14904 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _517_
timestamp 1
transform -1 0 16836 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _518_
timestamp 1
transform -1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _519_
timestamp 1
transform 1 0 14812 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _520_
timestamp 1
transform -1 0 14904 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _521_
timestamp 1
transform -1 0 16284 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _522_
timestamp 1
transform -1 0 12420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _523_
timestamp 1
transform 1 0 11592 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _524_
timestamp 1
transform -1 0 6808 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _525_
timestamp 1
transform 1 0 7176 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _526_
timestamp 1
transform -1 0 5612 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _527_
timestamp 1
transform 1 0 5796 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _528_
timestamp 1
transform 1 0 14168 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _529_
timestamp 1
transform -1 0 12052 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _530_
timestamp 1
transform 1 0 11592 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _531_
timestamp 1
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _532_
timestamp 1
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _533_
timestamp 1
transform -1 0 11408 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _534_
timestamp 1
transform 1 0 10856 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _535_
timestamp 1
transform -1 0 11040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _536_
timestamp 1
transform -1 0 10672 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _537_
timestamp 1
transform 1 0 9568 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _538_
timestamp 1
transform -1 0 12052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _539_
timestamp 1
transform 1 0 10580 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _540_
timestamp 1
transform 1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _541_
timestamp 1
transform 1 0 9660 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _542_
timestamp 1
transform -1 0 9384 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _543_
timestamp 1
transform -1 0 9660 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _544_
timestamp 1
transform -1 0 9752 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _545_
timestamp 1
transform -1 0 9660 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _546_
timestamp 1
transform 1 0 9016 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _547_
timestamp 1
transform -1 0 8372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _548_
timestamp 1
transform 1 0 8740 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _549_
timestamp 1
transform -1 0 8740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _550_
timestamp 1
transform 1 0 8188 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _551_
timestamp 1
transform 1 0 5336 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _552_
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _553_
timestamp 1
transform -1 0 6716 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _554_
timestamp 1
transform -1 0 7176 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _555_
timestamp 1
transform -1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _556_
timestamp 1
transform -1 0 7636 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _557_
timestamp 1
transform 1 0 7728 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _558_
timestamp 1
transform -1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _559_
timestamp 1
transform 1 0 7912 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_1  _560_
timestamp 1
transform 1 0 7176 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _561_
timestamp 1
transform 1 0 7544 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _562_
timestamp 1
transform -1 0 14720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _563_
timestamp 1
transform 1 0 12880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _564_
timestamp 1
transform 1 0 12512 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _565_
timestamp 1
transform -1 0 13616 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _566_
timestamp 1
transform -1 0 13800 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _567_
timestamp 1
transform -1 0 9568 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _568_
timestamp 1
transform -1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _569_
timestamp 1
transform -1 0 8648 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _570_
timestamp 1
transform 1 0 3772 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _571_
timestamp 1
transform 1 0 7636 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _572_
timestamp 1
transform 1 0 7544 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _573_
timestamp 1
transform 1 0 11040 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _574_
timestamp 1
transform 1 0 10948 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _575_
timestamp 1
transform -1 0 17388 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _576_
timestamp 1
transform 1 0 11868 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _577_
timestamp 1
transform 1 0 11776 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _578_
timestamp 1
transform -1 0 5704 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _579_
timestamp 1
transform 1 0 7820 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _580_
timestamp 1
transform 1 0 6992 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _581_
timestamp 1
transform -1 0 10488 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _582_
timestamp 1
transform 1 0 6532 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _583_
timestamp 1
transform 1 0 6992 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _584_
timestamp 1
transform -1 0 7820 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _585_
timestamp 1
transform 1 0 6716 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _586_
timestamp 1
transform 1 0 13708 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _587_
timestamp 1
transform 1 0 13248 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _588_
timestamp 1
transform -1 0 12236 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _589_
timestamp 1
transform 1 0 12420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _590_
timestamp 1
transform -1 0 13340 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _591_
timestamp 1
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _592_
timestamp 1
transform 1 0 14076 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _593_
timestamp 1
transform 1 0 13156 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _594_
timestamp 1
transform 1 0 13340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _595_
timestamp 1
transform -1 0 13984 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _596_
timestamp 1
transform 1 0 13432 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _597_
timestamp 1
transform 1 0 15640 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _598_
timestamp 1
transform 1 0 14628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _599_
timestamp 1
transform -1 0 14996 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _600_
timestamp 1
transform 1 0 14536 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _601_
timestamp 1
transform -1 0 13800 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _602_
timestamp 1
transform -1 0 14168 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _603_
timestamp 1
transform -1 0 16376 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _604_
timestamp 1
transform 1 0 14904 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _605_
timestamp 1
transform 1 0 12788 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _606_
timestamp 1
transform -1 0 14536 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _607_
timestamp 1
transform -1 0 11132 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _608_
timestamp 1
transform 1 0 9844 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _609_
timestamp 1
transform -1 0 11316 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _610_
timestamp 1
transform 1 0 14812 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _611_
timestamp 1
transform -1 0 14720 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _612_
timestamp 1
transform -1 0 14812 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _613_
timestamp 1
transform -1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _614_
timestamp 1
transform 1 0 9384 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _615_
timestamp 1
transform 1 0 8924 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _616_
timestamp 1
transform -1 0 10304 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _617_
timestamp 1
transform -1 0 11776 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _618_
timestamp 1
transform 1 0 12788 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _619_
timestamp 1
transform 1 0 13064 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o32ai_1  _620_
timestamp 1
transform -1 0 12972 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _621_
timestamp 1
transform -1 0 11316 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _622_
timestamp 1
transform -1 0 14628 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _623_
timestamp 1
transform 1 0 15364 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _624_
timestamp 1
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _625_
timestamp 1
transform -1 0 12236 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _626_
timestamp 1
transform 1 0 11132 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _627_
timestamp 1
transform 1 0 12328 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _628_
timestamp 1
transform -1 0 11868 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _629_
timestamp 1
transform 1 0 11960 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _630_
timestamp 1
transform 1 0 12052 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _631_
timestamp 1
transform -1 0 5520 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _632_
timestamp 1
transform -1 0 6624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _633_
timestamp 1
transform 1 0 7268 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _634_
timestamp 1
transform -1 0 3312 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _635_
timestamp 1
transform -1 0 1840 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _636_
timestamp 1
transform -1 0 5336 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _637_
timestamp 1
transform 1 0 3680 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _638_
timestamp 1
transform 1 0 4232 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _639_
timestamp 1
transform 1 0 3588 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _640_
timestamp 1
transform 1 0 5428 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _641_
timestamp 1
transform -1 0 11592 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _642_
timestamp 1
transform 1 0 5704 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _643_
timestamp 1
transform 1 0 4784 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _644_
timestamp 1
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _645_
timestamp 1
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _646_
timestamp 1
transform -1 0 5520 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _647_
timestamp 1
transform -1 0 3496 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _648_
timestamp 1
transform 1 0 2576 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _649_
timestamp 1
transform 1 0 2300 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _650_
timestamp 1
transform -1 0 2760 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _651_
timestamp 1
transform 1 0 1472 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _652_
timestamp 1
transform 1 0 12788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _653_
timestamp 1
transform -1 0 12604 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _654_
timestamp 1
transform -1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _655_
timestamp 1
transform 1 0 12236 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _656_
timestamp 1
transform -1 0 12236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _657_
timestamp 1
transform 1 0 11776 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _658_
timestamp 1
transform 1 0 12512 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _659_
timestamp 1
transform 1 0 12420 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _660_
timestamp 1
transform 1 0 12236 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _661_
timestamp 1
transform 1 0 15640 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _662_
timestamp 1
transform 1 0 14904 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _663_
timestamp 1
transform -1 0 15640 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _664_
timestamp 1
transform -1 0 13892 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _665_
timestamp 1
transform -1 0 14260 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _666_
timestamp 1
transform -1 0 12512 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _667_
timestamp 1
transform -1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _668_
timestamp 1
transform 1 0 13064 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _669_
timestamp 1
transform 1 0 12972 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_1  _670_
timestamp 1
transform 1 0 12696 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _671_
timestamp 1
transform -1 0 8188 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _672_
timestamp 1
transform 1 0 7084 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _673_
timestamp 1
transform 1 0 6992 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _674_
timestamp 1
transform 1 0 5060 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _675_
timestamp 1
transform -1 0 7176 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _676_
timestamp 1
transform 1 0 6440 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _677_
timestamp 1
transform 1 0 5244 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _678_
timestamp 1
transform -1 0 10856 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _679_
timestamp 1
transform 1 0 9476 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _680_
timestamp 1
transform 1 0 2392 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _681_
timestamp 1
transform 1 0 2760 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _682_
timestamp 1
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _683_
timestamp 1
transform 1 0 3864 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _684_
timestamp 1
transform -1 0 4600 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _685_
timestamp 1
transform 1 0 3772 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _686_
timestamp 1
transform -1 0 6256 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _687_
timestamp 1
transform 1 0 3956 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _688_
timestamp 1
transform 1 0 2300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _689_
timestamp 1
transform 1 0 2116 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _690_
timestamp 1
transform -1 0 2116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _691_
timestamp 1
transform -1 0 4508 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _692_
timestamp 1
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _693_
timestamp 1
transform 1 0 3036 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _694_
timestamp 1
transform -1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _695_
timestamp 1
transform 1 0 3864 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _696_
timestamp 1
transform 1 0 5428 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _697_
timestamp 1
transform 1 0 4232 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _698_
timestamp 1
transform 1 0 6348 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _699_
timestamp 1
transform -1 0 7084 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_1  _700_
timestamp 1
transform -1 0 6624 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _701_
timestamp 1
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _702_
timestamp 1
transform 1 0 2484 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _703_
timestamp 1
transform -1 0 11316 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _704_
timestamp 1
transform 1 0 2576 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _705_
timestamp 1
transform 1 0 4324 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _706_
timestamp 1
transform 1 0 3772 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _707_
timestamp 1
transform 1 0 2300 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _708_
timestamp 1
transform 1 0 2944 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _709_
timestamp 1
transform -1 0 3404 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _710_
timestamp 1
transform -1 0 2852 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _711_
timestamp 1
transform -1 0 2208 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _712_
timestamp 1
transform 1 0 10672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _713_
timestamp 1
transform 1 0 10396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _714_
timestamp 1
transform 1 0 9016 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _715_
timestamp 1
transform 1 0 6348 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _716_
timestamp 1
transform 1 0 10856 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _717_
timestamp 1
transform 1 0 11684 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _718_
timestamp 1
transform -1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _719_
timestamp 1
transform 1 0 8924 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _720_
timestamp 1
transform 1 0 8832 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _721_
timestamp 1
transform 1 0 9752 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _722_
timestamp 1
transform 1 0 9660 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _723_
timestamp 1
transform 1 0 9384 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _724_
timestamp 1
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _725_
timestamp 1
transform -1 0 9752 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _726_
timestamp 1
transform 1 0 9752 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _727_
timestamp 1
transform 1 0 10028 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _728_
timestamp 1
transform -1 0 9108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _729_
timestamp 1
transform -1 0 9200 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _730_
timestamp 1
transform 1 0 6900 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _731_
timestamp 1
transform 1 0 5244 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _732_
timestamp 1
transform -1 0 5888 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _733_
timestamp 1
transform 1 0 7728 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _734_
timestamp 1
transform 1 0 12420 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _735_
timestamp 1
transform -1 0 12972 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _736_
timestamp 1
transform 1 0 12972 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _737_
timestamp 1
transform 1 0 7636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _738_
timestamp 1
transform 1 0 5520 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _739_
timestamp 1
transform 1 0 7452 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _740_
timestamp 1
transform -1 0 4600 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _741_
timestamp 1
transform 1 0 3312 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _742_
timestamp 1
transform 1 0 2852 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _743_
timestamp 1
transform -1 0 4968 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _744_
timestamp 1
transform -1 0 4416 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _745_
timestamp 1
transform 1 0 3864 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _746_
timestamp 1
transform 1 0 3220 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _747_
timestamp 1
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _748_
timestamp 1
transform -1 0 12144 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _749_
timestamp 1
transform 1 0 10764 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _750_
timestamp 1
transform -1 0 9844 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _751_
timestamp 1
transform -1 0 11132 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _752_
timestamp 1
transform 1 0 15272 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _753_
timestamp 1
transform 1 0 15456 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _754_
timestamp 1
transform -1 0 15088 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _755_
timestamp 1
transform -1 0 15456 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _756_
timestamp 1
transform 1 0 15088 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _757_
timestamp 1
transform -1 0 15548 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _758_
timestamp 1
transform -1 0 17296 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _759_
timestamp 1
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _760_
timestamp 1
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _761_
timestamp 1
transform -1 0 16192 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _762_
timestamp 1
transform 1 0 4508 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _763_
timestamp 1
transform -1 0 6164 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _764_
timestamp 1
transform 1 0 5152 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _765_
timestamp 1
transform -1 0 4508 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _766_
timestamp 1
transform 1 0 6624 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _767_
timestamp 1
transform -1 0 8188 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _768_
timestamp 1
transform -1 0 7176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _769_
timestamp 1
transform 1 0 7728 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _770_
timestamp 1
transform 1 0 6900 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _771_
timestamp 1
transform -1 0 11316 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _772_
timestamp 1
transform -1 0 8832 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _773_
timestamp 1
transform 1 0 7544 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _774_
timestamp 1
transform 1 0 9844 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _775_
timestamp 1
transform 1 0 10304 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _776_
timestamp 1
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _777_
timestamp 1
transform -1 0 11316 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a32oi_2  _778_
timestamp 1
transform 1 0 8648 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _779_
timestamp 1
transform -1 0 10120 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _780_
timestamp 1
transform 1 0 9200 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _781_
timestamp 1
transform -1 0 9200 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _782_
timestamp 1
transform 1 0 9660 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _783_
timestamp 1
transform -1 0 13156 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _784_
timestamp 1
transform 1 0 13616 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _785_
timestamp 1
transform 1 0 13616 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _786_
timestamp 1
transform 1 0 12788 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _787_
timestamp 1
transform 1 0 13800 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _788_
timestamp 1
transform -1 0 13800 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _789_
timestamp 1
transform 1 0 13432 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _790_
timestamp 1
transform 1 0 12972 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _791_
timestamp 1
transform -1 0 17664 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _792_
timestamp 1
transform 1 0 17664 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _793_
timestamp 1
transform -1 0 16928 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _794_
timestamp 1
transform -1 0 16192 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _795_
timestamp 1
transform -1 0 16652 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _796_
timestamp 1
transform -1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _797_
timestamp 1
transform -1 0 16836 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _798_
timestamp 1
transform -1 0 17756 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _799_
timestamp 1
transform 1 0 16192 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _800_
timestamp 1
transform -1 0 18124 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _801_
timestamp 1
transform 1 0 15272 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _802_
timestamp 1
transform 1 0 14076 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _803_
timestamp 1
transform 1 0 13984 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _804_
timestamp 1
transform 1 0 14444 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _805_
timestamp 1
transform 1 0 14444 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform -1 0 16560 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1
transform 1 0 16284 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1
transform -1 0 16560 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout19
timestamp 1
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout20
timestamp 1
transform 1 0 14352 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout21
timestamp 1
transform -1 0 10212 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 1
transform 1 0 4968 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1
transform -1 0 17388 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 1
transform 1 0 15824 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout25
timestamp 1
transform 1 0 16744 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout26
timestamp 1
transform -1 0 14444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout27
timestamp 1
transform -1 0 10120 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 1
transform 1 0 15824 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1
transform -1 0 13892 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout30
timestamp 1
transform 1 0 14812 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1
transform 1 0 14904 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout32
timestamp 1
transform -1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout33
timestamp 1
transform -1 0 16376 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout34
timestamp 1
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 1
transform -1 0 9936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout36
timestamp 1
transform -1 0 7728 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 1
transform 1 0 15180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout38
timestamp 1
transform -1 0 15916 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout39
timestamp 1
transform 1 0 16652 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp 1
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 1
transform -1 0 8648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp 1
transform 1 0 15088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout43
timestamp 1
transform 1 0 13248 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout44
timestamp 1
transform -1 0 14996 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout45
timestamp 1
transform 1 0 4876 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout46
timestamp 1
transform -1 0 7636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp 1
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout48
timestamp 1
transform -1 0 6164 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout49
timestamp 1
transform -1 0 8832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout50
timestamp 1
transform -1 0 13248 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout51
timestamp 1
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout52
timestamp 1
transform 1 0 12696 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout53
timestamp 1
transform -1 0 16008 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout54
timestamp 1
transform -1 0 16376 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout55
timestamp 1
transform 1 0 5888 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout56
timestamp 1
transform -1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout57
timestamp 1
transform 1 0 9292 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout58
timestamp 1
transform -1 0 10212 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout59
timestamp 1
transform 1 0 14720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp 1
transform 1 0 17020 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout61
timestamp 1
transform 1 0 17020 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout62
timestamp 1
transform -1 0 6440 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout63
timestamp 1
transform -1 0 6256 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout64
timestamp 1
transform -1 0 9844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout65
timestamp 1
transform 1 0 17572 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout66
timestamp 1
transform 1 0 16744 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout67
timestamp 1
transform -1 0 5888 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout68
timestamp 1
transform -1 0 4876 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  fanout69
timestamp 1
transform -1 0 9108 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout70
timestamp 1
transform -1 0 10028 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout71
timestamp 1
transform -1 0 17296 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout72
timestamp 1
transform 1 0 15824 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63
timestamp 1636968456
transform 1 0 6900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75
timestamp 1
transform 1 0 8004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98
timestamp 1636968456
transform 1 0 10120 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125
timestamp 1
transform 1 0 12604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_133
timestamp 1
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636968456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 1
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_85
timestamp 1
transform 1 0 8924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_103
timestamp 1
transform 1 0 10580 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_113
timestamp 1
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_119
timestamp 1
transform 1 0 12052 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_123
timestamp 1
transform 1 0 12420 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_136
timestamp 1636968456
transform 1 0 13616 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_148
timestamp 1636968456
transform 1 0 14720 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_160
timestamp 1
transform 1 0 15824 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_19
timestamp 1
transform 1 0 2852 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp 1
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_50
timestamp 1
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_75
timestamp 1
transform 1 0 8004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_100
timestamp 1
transform 1 0 10304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_111
timestamp 1
transform 1 0 11316 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_125
timestamp 1
transform 1 0 12604 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_146
timestamp 1
transform 1 0 14536 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp 1
transform 1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_156
timestamp 1636968456
transform 1 0 15456 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_168
timestamp 1636968456
transform 1 0 16560 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_184
timestamp 1
transform 1 0 18032 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1
transform 1 0 2484 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_45
timestamp 1
transform 1 0 5244 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_69
timestamp 1
transform 1 0 7452 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_99
timestamp 1
transform 1 0 10212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 1
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_121
timestamp 1
transform 1 0 12236 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_129
timestamp 1
transform 1 0 12972 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_138
timestamp 1
transform 1 0 13800 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_146
timestamp 1
transform 1 0 14536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_178
timestamp 1
transform 1 0 17480 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_184
timestamp 1
transform 1 0 18032 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_19
timestamp 1
transform 1 0 2852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_54
timestamp 1
transform 1 0 6072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_73
timestamp 1
transform 1 0 7820 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636968456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_114
timestamp 1
transform 1 0 11592 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_121
timestamp 1
transform 1 0 12236 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_129
timestamp 1
transform 1 0 12972 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_145
timestamp 1
transform 1 0 14444 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_151
timestamp 1
transform 1 0 14996 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_166
timestamp 1636968456
transform 1 0 16376 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_178
timestamp 1
transform 1 0 17480 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_184
timestamp 1
transform 1 0 18032 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636968456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636968456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1
transform 1 0 3588 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_36
timestamp 1636968456
transform 1 0 4416 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_48
timestamp 1
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636968456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_81
timestamp 1
transform 1 0 8556 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_88
timestamp 1
transform 1 0 9200 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_96
timestamp 1
transform 1 0 9936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp 1
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_113
timestamp 1
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_119
timestamp 1
transform 1 0 12052 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_146
timestamp 1
transform 1 0 14536 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_150
timestamp 1
transform 1 0 14904 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636968456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7
timestamp 1636968456
transform 1 0 1748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_19
timestamp 1
transform 1 0 2852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_37
timestamp 1
transform 1 0 4508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_46
timestamp 1
transform 1 0 5336 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_55
timestamp 1
transform 1 0 6164 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_94
timestamp 1
transform 1 0 9752 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_111
timestamp 1
transform 1 0 11316 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_122
timestamp 1
transform 1 0 12328 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_126
timestamp 1
transform 1 0 12696 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_130
timestamp 1
transform 1 0 13064 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp 1
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_157
timestamp 1
transform 1 0 15548 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_176
timestamp 1
transform 1 0 17296 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_184
timestamp 1
transform 1 0 18032 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636968456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp 1
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_42
timestamp 1
transform 1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_52
timestamp 1
transform 1 0 5888 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_61
timestamp 1
transform 1 0 6716 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_68
timestamp 1
transform 1 0 7360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_79
timestamp 1
transform 1 0 8372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_101
timestamp 1
transform 1 0 10396 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_136
timestamp 1
transform 1 0 13616 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_156
timestamp 1
transform 1 0 15456 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_182
timestamp 1
transform 1 0 17848 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636968456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_58
timestamp 1
transform 1 0 6440 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_74
timestamp 1
transform 1 0 7912 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636968456
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636968456
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_109
timestamp 1
transform 1 0 11132 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_120
timestamp 1636968456
transform 1 0 12144 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_132
timestamp 1
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_141
timestamp 1
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_157
timestamp 1
transform 1 0 15548 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_165
timestamp 1
transform 1 0 16284 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_172
timestamp 1636968456
transform 1 0 16928 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_184
timestamp 1
transform 1 0 18032 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636968456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_22
timestamp 1
transform 1 0 3128 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_38
timestamp 1
transform 1 0 4600 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_44
timestamp 1
transform 1 0 5152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_65
timestamp 1
transform 1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_75
timestamp 1
transform 1 0 8004 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_83
timestamp 1
transform 1 0 8740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_94
timestamp 1
transform 1 0 9752 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_119
timestamp 1
transform 1 0 12052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_142
timestamp 1
transform 1 0 14168 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_150
timestamp 1
transform 1 0 14904 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_169
timestamp 1
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_176
timestamp 1
transform 1 0 17296 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_184
timestamp 1
transform 1 0 18032 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636968456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_15
timestamp 1
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_22
timestamp 1
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_35
timestamp 1
transform 1 0 4324 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_39
timestamp 1
transform 1 0 4692 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_71
timestamp 1636968456
transform 1 0 7636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_101
timestamp 1
transform 1 0 10396 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_105
timestamp 1
transform 1 0 10764 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_122
timestamp 1
transform 1 0 12328 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_130
timestamp 1
transform 1 0 13064 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_149
timestamp 1
transform 1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_157
timestamp 1
transform 1 0 15548 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_162
timestamp 1636968456
transform 1 0 16008 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_174
timestamp 1
transform 1 0 17112 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_180
timestamp 1
transform 1 0 17664 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636968456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636968456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_31
timestamp 1
transform 1 0 3956 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_37
timestamp 1
transform 1 0 4508 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_45
timestamp 1
transform 1 0 5244 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_85
timestamp 1
transform 1 0 8924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_102
timestamp 1
transform 1 0 10488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_121
timestamp 1
transform 1 0 12236 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_174
timestamp 1
transform 1 0 17112 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_182
timestamp 1
transform 1 0 17848 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_7
timestamp 1
transform 1 0 1748 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_19
timestamp 1
transform 1 0 2852 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_38
timestamp 1
transform 1 0 4600 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_45
timestamp 1
transform 1 0 5244 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_53
timestamp 1
transform 1 0 5980 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_60
timestamp 1
transform 1 0 6624 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_66
timestamp 1
transform 1 0 7176 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_71
timestamp 1
transform 1 0 7636 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_85
timestamp 1
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_99
timestamp 1636968456
transform 1 0 10212 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_111
timestamp 1
transform 1 0 11316 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_122
timestamp 1636968456
transform 1 0 12328 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_166
timestamp 1
transform 1 0 16376 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_178
timestamp 1
transform 1 0 17480 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_184
timestamp 1
transform 1 0 18032 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_12
timestamp 1
transform 1 0 2208 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_30
timestamp 1
transform 1 0 3864 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_75
timestamp 1636968456
transform 1 0 8004 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_87
timestamp 1
transform 1 0 9108 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_93
timestamp 1
transform 1 0 9660 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_99
timestamp 1636968456
transform 1 0 10212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 1
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1
transform 1 0 13248 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_136
timestamp 1
transform 1 0 13616 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_152
timestamp 1
transform 1 0 15088 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_160
timestamp 1
transform 1 0 15824 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636968456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_36
timestamp 1
transform 1 0 4416 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_58
timestamp 1
transform 1 0 6440 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_72
timestamp 1
transform 1 0 7728 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_80
timestamp 1
transform 1 0 8464 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_98
timestamp 1
transform 1 0 10120 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_141
timestamp 1
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1
transform 1 0 14812 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_153
timestamp 1
transform 1 0 15180 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_159
timestamp 1
transform 1 0 15732 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_177
timestamp 1
transform 1 0 17388 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636968456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_15
timestamp 1
transform 1 0 2484 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_24
timestamp 1
transform 1 0 3312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_57
timestamp 1
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_66
timestamp 1636968456
transform 1 0 7176 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_78
timestamp 1
transform 1 0 8280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_82
timestamp 1
transform 1 0 8648 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_93
timestamp 1
transform 1 0 9660 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_102
timestamp 1
transform 1 0 10488 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_106
timestamp 1
transform 1 0 10856 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_129
timestamp 1
transform 1 0 12972 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_137
timestamp 1
transform 1 0 13708 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_148
timestamp 1
transform 1 0 14720 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_161
timestamp 1
transform 1 0 15916 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_177
timestamp 1
transform 1 0 17388 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_35
timestamp 1
transform 1 0 4324 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_41
timestamp 1
transform 1 0 4876 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_57
timestamp 1
transform 1 0 6348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_65
timestamp 1
transform 1 0 7084 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_69
timestamp 1
transform 1 0 7452 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_89
timestamp 1
transform 1 0 9292 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_104
timestamp 1
transform 1 0 10672 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_123
timestamp 1
transform 1 0 12420 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_131
timestamp 1
transform 1 0 13156 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_184
timestamp 1
transform 1 0 18032 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_11
timestamp 1
transform 1 0 2116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_23
timestamp 1
transform 1 0 3220 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp 1
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_36
timestamp 1636968456
transform 1 0 4416 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_48
timestamp 1
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_57
timestamp 1
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_80
timestamp 1
transform 1 0 8464 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_88
timestamp 1
transform 1 0 9200 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_101
timestamp 1
transform 1 0 10396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_126
timestamp 1
transform 1 0 12696 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_131
timestamp 1
transform 1 0 13156 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1
transform 1 0 13892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1
transform 1 0 14352 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_148
timestamp 1
transform 1 0 14720 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_154
timestamp 1636968456
transform 1 0 15272 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_174
timestamp 1
transform 1 0 17112 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_182
timestamp 1
transform 1 0 17848 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_11
timestamp 1
transform 1 0 2116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_22
timestamp 1
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_42
timestamp 1
transform 1 0 4968 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_52
timestamp 1
transform 1 0 5888 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_58
timestamp 1
transform 1 0 6440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_90
timestamp 1
transform 1 0 9384 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_95
timestamp 1636968456
transform 1 0 9844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_107
timestamp 1
transform 1 0 10948 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_120
timestamp 1
transform 1 0 12144 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_124
timestamp 1
transform 1 0 12512 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_141
timestamp 1
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_151
timestamp 1
transform 1 0 14996 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_159
timestamp 1
transform 1 0 15732 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_181
timestamp 1
transform 1 0 17756 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_13
timestamp 1
transform 1 0 2300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_22
timestamp 1
transform 1 0 3128 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_26
timestamp 1
transform 1 0 3496 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_44
timestamp 1
transform 1 0 5152 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_65
timestamp 1636968456
transform 1 0 7084 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_77
timestamp 1
transform 1 0 8188 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_88
timestamp 1
transform 1 0 9200 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_98
timestamp 1
transform 1 0 10120 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_121
timestamp 1
transform 1 0 12236 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_129
timestamp 1
transform 1 0 12972 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_145
timestamp 1
transform 1 0 14444 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_173
timestamp 1
transform 1 0 17020 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_183
timestamp 1
transform 1 0 17940 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_34
timestamp 1
transform 1 0 4232 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_42
timestamp 1
transform 1 0 4968 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_48
timestamp 1636968456
transform 1 0 5520 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_60
timestamp 1
transform 1 0 6624 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_64
timestamp 1
transform 1 0 6992 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_72
timestamp 1
transform 1 0 7728 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_80
timestamp 1
transform 1 0 8464 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_100
timestamp 1
transform 1 0 10304 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_104
timestamp 1
transform 1 0 10672 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_112
timestamp 1636968456
transform 1 0 11408 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_124
timestamp 1
transform 1 0 12512 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_149
timestamp 1
transform 1 0 14812 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_156
timestamp 1
transform 1 0 15456 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_164
timestamp 1
transform 1 0 16192 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_7
timestamp 1
transform 1 0 1748 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_24
timestamp 1
transform 1 0 3312 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_34
timestamp 1
transform 1 0 4232 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_42
timestamp 1
transform 1 0 4968 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_47
timestamp 1
transform 1 0 5428 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_57
timestamp 1
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_71
timestamp 1
transform 1 0 7636 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_88
timestamp 1
transform 1 0 9200 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_99
timestamp 1
transform 1 0 10212 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_105
timestamp 1
transform 1 0 10764 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_121
timestamp 1636968456
transform 1 0 12236 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_133
timestamp 1
transform 1 0 13340 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_139
timestamp 1
transform 1 0 13892 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1
transform 1 0 17572 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_7
timestamp 1
transform 1 0 1748 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_17
timestamp 1
transform 1 0 2668 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_46
timestamp 1
transform 1 0 5336 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_74
timestamp 1
transform 1 0 7912 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_80
timestamp 1
transform 1 0 8464 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_100
timestamp 1
transform 1 0 10304 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_108
timestamp 1
transform 1 0 11040 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_117
timestamp 1
transform 1 0 11868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_121
timestamp 1
transform 1 0 12236 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_129
timestamp 1
transform 1 0 12972 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_25
timestamp 1
transform 1 0 3404 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_35
timestamp 1636968456
transform 1 0 4324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_47
timestamp 1
transform 1 0 5428 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_57
timestamp 1
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_63
timestamp 1
transform 1 0 6900 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_77
timestamp 1
transform 1 0 8188 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_83
timestamp 1
transform 1 0 8740 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_87
timestamp 1
transform 1 0 9108 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_97
timestamp 1
transform 1 0 10028 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1
transform 1 0 12144 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_137
timestamp 1
transform 1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_145
timestamp 1
transform 1 0 14444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_177
timestamp 1
transform 1 0 17388 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_11
timestamp 1
transform 1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_29
timestamp 1
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_38
timestamp 1
transform 1 0 4600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_61
timestamp 1
transform 1 0 6716 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_69
timestamp 1
transform 1 0 7452 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_100
timestamp 1636968456
transform 1 0 10304 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_112
timestamp 1636968456
transform 1 0 11408 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_124
timestamp 1
transform 1 0 12512 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_130
timestamp 1
transform 1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_149
timestamp 1
transform 1 0 14812 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_182
timestamp 1
transform 1 0 17848 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636968456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_15
timestamp 1
transform 1 0 2484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_39
timestamp 1
transform 1 0 4692 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_73
timestamp 1
transform 1 0 7820 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_79
timestamp 1
transform 1 0 8372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_87
timestamp 1
transform 1 0 9108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_100
timestamp 1
transform 1 0 10304 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_172
timestamp 1
transform 1 0 16928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_177
timestamp 1
transform 1 0 17388 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636968456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_15
timestamp 1
transform 1 0 2484 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_29
timestamp 1
transform 1 0 3772 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_55
timestamp 1
transform 1 0 6164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_79
timestamp 1
transform 1 0 8372 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_111
timestamp 1636968456
transform 1 0 11316 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_123
timestamp 1
transform 1 0 12420 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_127
timestamp 1
transform 1 0 12788 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_131
timestamp 1
transform 1 0 13156 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_169
timestamp 1636968456
transform 1 0 16652 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_181
timestamp 1
transform 1 0 17756 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636968456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1636968456
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_27
timestamp 1
transform 1 0 3588 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_34
timestamp 1
transform 1 0 4232 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_42
timestamp 1
transform 1 0 4968 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_66
timestamp 1
transform 1 0 7176 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_76
timestamp 1
transform 1 0 8096 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_102
timestamp 1
transform 1 0 10488 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_122
timestamp 1
transform 1 0 12328 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_130
timestamp 1
transform 1 0 13064 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_143
timestamp 1
transform 1 0 14260 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_147
timestamp 1
transform 1 0 14628 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_175
timestamp 1
transform 1 0 17204 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_183
timestamp 1
transform 1 0 17940 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636968456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_15
timestamp 1
transform 1 0 2484 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636968456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636968456
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1636968456
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1636968456
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 1
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_98
timestamp 1
transform 1 0 10120 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_105
timestamp 1
transform 1 0 10764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_117
timestamp 1
transform 1 0 11868 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_123
timestamp 1
transform 1 0 12420 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_171
timestamp 1636968456
transform 1 0 16836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_183
timestamp 1
transform 1 0 17940 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636968456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636968456
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1636968456
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1636968456
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636968456
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_69
timestamp 1
transform 1 0 7452 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_92
timestamp 1
transform 1 0 9568 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_98
timestamp 1
transform 1 0 10120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_123
timestamp 1
transform 1 0 12420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_139
timestamp 1
transform 1 0 13892 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1636968456
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_181
timestamp 1
transform 1 0 17756 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636968456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636968456
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1636968456
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1636968456
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_53
timestamp 1
transform 1 0 5980 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_57
timestamp 1636968456
transform 1 0 6348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_69
timestamp 1
transform 1 0 7452 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_77
timestamp 1
transform 1 0 8188 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_85
timestamp 1
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_93
timestamp 1
transform 1 0 9660 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_98
timestamp 1
transform 1 0 10120 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_105
timestamp 1
transform 1 0 10764 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_113
timestamp 1636968456
transform 1 0 11500 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_125
timestamp 1
transform 1 0 12604 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_131
timestamp 1
transform 1 0 13156 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_165
timestamp 1
transform 1 0 16284 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_169
timestamp 1636968456
transform 1 0 16652 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1
transform -1 0 18124 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  max_cap18
timestamp 1
transform 1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output2
timestamp 1
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1
transform 1 0 17756 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1
transform 1 0 7820 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1
transform 1 0 11040 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1
transform 1 0 9752 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1
transform 1 0 10396 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1
transform -1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1
transform 1 0 17756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_31
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 18400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_32
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 18400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_33
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_34
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 18400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_35
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 18400 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_36
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 18400 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_37
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 18400 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_38
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 18400 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_39
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 18400 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_40
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 18400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_41
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 18400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_42
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 18400 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_43
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 18400 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_44
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 18400 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_45
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 18400 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_46
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 18400 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_47
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 18400 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_48
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 18400 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_49
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 18400 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_50
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 18400 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_51
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 18400 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_52
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 18400 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_53
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 18400 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_54
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 18400 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_55
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 18400 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_56
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 18400 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_57
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 18400 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_58
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 18400 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_59
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 18400 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_60
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 18400 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_61
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 18400 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_64
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_65
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_66
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_67
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_68
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_69
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_70
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_71
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_72
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_73
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_74
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_75
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_76
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_77
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_78
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_79
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_80
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_81
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_82
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_83
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_84
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_85
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_87
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_88
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_92
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_93
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_95
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_96
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_97
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_98
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_99
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_100
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_101
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_102
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_103
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_104
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_105
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_106
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_107
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_108
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_109
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_110
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_111
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_112
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_113
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_114
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_115
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_116
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_117
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_118
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_119
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_120
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_121
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_122
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_123
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_124
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_125
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_126
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_127
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_128
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_129
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_130
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_131
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_132
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_133
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_134
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_135
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_136
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_137
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_138
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_139
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_140
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_141
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_142
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_143
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_144
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_145
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_146
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_147
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_148
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_149
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_150
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_151
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_152
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_153
timestamp 1
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_154
timestamp 1
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_155
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_156
timestamp 1
transform 1 0 6256 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_157
timestamp 1
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_158
timestamp 1
transform 1 0 11408 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_159
timestamp 1
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_160
timestamp 1
transform 1 0 16560 0 1 18496
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 18760 13608 19560 13728 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 18760 14968 19560 15088 0 FreeSans 480 0 0 0 rst
port 3 nsew signal input
flabel metal2 s 8390 20904 8446 21704 0 FreeSans 224 90 0 0 sine_out[0]
port 4 nsew signal output
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 sine_out[10]
port 5 nsew signal output
flabel metal3 s 18760 14288 19560 14408 0 FreeSans 480 0 0 0 sine_out[11]
port 6 nsew signal output
flabel metal2 s 7746 20904 7802 21704 0 FreeSans 224 90 0 0 sine_out[12]
port 7 nsew signal output
flabel metal2 s 10966 20904 11022 21704 0 FreeSans 224 90 0 0 sine_out[13]
port 8 nsew signal output
flabel metal2 s 9678 20904 9734 21704 0 FreeSans 224 90 0 0 sine_out[14]
port 9 nsew signal output
flabel metal2 s 10322 20904 10378 21704 0 FreeSans 224 90 0 0 sine_out[15]
port 10 nsew signal output
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 sine_out[1]
port 11 nsew signal output
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 sine_out[2]
port 12 nsew signal output
flabel metal3 s 18760 7488 19560 7608 0 FreeSans 480 0 0 0 sine_out[3]
port 13 nsew signal output
flabel metal2 s 12898 20904 12954 21704 0 FreeSans 224 90 0 0 sine_out[4]
port 14 nsew signal output
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 sine_out[5]
port 15 nsew signal output
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 sine_out[6]
port 16 nsew signal output
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 sine_out[7]
port 17 nsew signal output
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 sine_out[8]
port 18 nsew signal output
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 sine_out[9]
port 19 nsew signal output
rlabel metal1 9752 18496 9752 18496 0 VGND
rlabel metal1 9752 19040 9752 19040 0 VPWR
rlabel metal1 16790 10778 16790 10778 0 _000_
rlabel metal1 16054 13158 16054 13158 0 _001_
rlabel metal2 17526 14178 17526 14178 0 _002_
rlabel metal1 15318 15402 15318 15402 0 _003_
rlabel metal1 14214 16014 14214 16014 0 _004_
rlabel metal1 13386 18360 13386 18360 0 _005_
rlabel metal1 14306 17714 14306 17714 0 _006_
rlabel metal1 14122 17850 14122 17850 0 _007_
rlabel metal1 16836 12682 16836 12682 0 _008_
rlabel metal2 17526 11832 17526 11832 0 _009_
rlabel metal1 17572 12954 17572 12954 0 _010_
rlabel metal2 16698 15674 16698 15674 0 _011_
rlabel metal1 15831 16150 15831 16150 0 _012_
rlabel metal2 16514 17442 16514 17442 0 _013_
rlabel metal2 15870 17850 15870 17850 0 _014_
rlabel metal2 16698 18258 16698 18258 0 _015_
rlabel metal1 10212 13362 10212 13362 0 _016_
rlabel metal1 9706 13328 9706 13328 0 _017_
rlabel via3 3059 12580 3059 12580 0 _018_
rlabel metal1 9154 4046 9154 4046 0 _019_
rlabel metal2 9246 5695 9246 5695 0 _020_
rlabel metal1 15226 6800 15226 6800 0 _021_
rlabel metal2 12650 10370 12650 10370 0 _022_
rlabel metal1 12512 12206 12512 12206 0 _023_
rlabel metal1 9016 10098 9016 10098 0 _024_
rlabel metal2 6026 5916 6026 5916 0 _025_
rlabel metal1 5290 8466 5290 8466 0 _026_
rlabel metal2 9614 13634 9614 13634 0 _027_
rlabel metal2 12466 7684 12466 7684 0 _028_
rlabel metal2 12558 10285 12558 10285 0 _029_
rlabel metal1 9476 13362 9476 13362 0 _030_
rlabel metal1 11178 5304 11178 5304 0 _031_
rlabel metal1 9522 6256 9522 6256 0 _032_
rlabel via2 9522 10251 9522 10251 0 _033_
rlabel metal1 8510 13498 8510 13498 0 _034_
rlabel via2 9338 15419 9338 15419 0 _035_
rlabel metal2 11546 6018 11546 6018 0 _036_
rlabel metal1 14444 5610 14444 5610 0 _037_
rlabel metal2 8602 12087 8602 12087 0 _038_
rlabel metal2 7360 8398 7360 8398 0 _039_
rlabel metal2 8050 11968 8050 11968 0 _040_
rlabel metal1 5658 4624 5658 4624 0 _041_
rlabel metal2 15226 9214 15226 9214 0 _042_
rlabel metal1 7590 13838 7590 13838 0 _043_
rlabel via1 6578 13838 6578 13838 0 _044_
rlabel metal2 14674 9027 14674 9027 0 _045_
rlabel metal1 3036 11866 3036 11866 0 _046_
rlabel metal2 3634 8806 3634 8806 0 _047_
rlabel metal1 4554 13498 4554 13498 0 _048_
rlabel metal1 9062 13430 9062 13430 0 _049_
rlabel metal2 7130 13702 7130 13702 0 _050_
rlabel via2 12834 15045 12834 15045 0 _051_
rlabel metal2 7498 15453 7498 15453 0 _052_
rlabel metal1 7774 13906 7774 13906 0 _053_
rlabel metal1 9522 11560 9522 11560 0 _054_
rlabel metal1 9982 7514 9982 7514 0 _055_
rlabel metal1 16238 8398 16238 8398 0 _056_
rlabel metal1 9936 9554 9936 9554 0 _057_
rlabel metal1 4508 12750 4508 12750 0 _058_
rlabel metal1 4232 13906 4232 13906 0 _059_
rlabel metal2 12558 13401 12558 13401 0 _060_
rlabel metal2 10074 8602 10074 8602 0 _061_
rlabel metal1 7682 7310 7682 7310 0 _062_
rlabel metal1 6670 12784 6670 12784 0 _063_
rlabel metal1 11730 16116 11730 16116 0 _064_
rlabel viali 9246 11119 9246 11119 0 _065_
rlabel metal1 6624 4590 6624 4590 0 _066_
rlabel via2 14398 12189 14398 12189 0 _067_
rlabel metal1 6072 7514 6072 7514 0 _068_
rlabel metal2 11178 10030 11178 10030 0 _069_
rlabel metal1 4508 7854 4508 7854 0 _070_
rlabel metal1 5888 7922 5888 7922 0 _071_
rlabel metal1 6233 10642 6233 10642 0 _072_
rlabel metal1 5934 7786 5934 7786 0 _073_
rlabel metal1 5842 10710 5842 10710 0 _074_
rlabel metal1 7084 6426 7084 6426 0 _075_
rlabel metal1 7728 13158 7728 13158 0 _076_
rlabel metal1 7314 6732 7314 6732 0 _077_
rlabel metal2 7774 7174 7774 7174 0 _078_
rlabel metal2 7682 7667 7682 7667 0 _079_
rlabel metal1 8648 7242 8648 7242 0 _080_
rlabel metal1 14858 6358 14858 6358 0 _081_
rlabel metal2 15778 10914 15778 10914 0 _082_
rlabel metal1 16054 8058 16054 8058 0 _083_
rlabel metal2 14582 6460 14582 6460 0 _084_
rlabel metal2 14398 6766 14398 6766 0 _085_
rlabel metal1 15594 7412 15594 7412 0 _086_
rlabel metal1 12190 3162 12190 3162 0 _087_
rlabel metal1 11408 7922 11408 7922 0 _088_
rlabel metal1 6348 15878 6348 15878 0 _089_
rlabel metal1 7682 15402 7682 15402 0 _090_
rlabel metal3 5727 9452 5727 9452 0 _091_
rlabel metal2 6210 7378 6210 7378 0 _092_
rlabel metal2 11822 7106 11822 7106 0 _093_
rlabel metal1 11638 7514 11638 7514 0 _094_
rlabel metal2 11178 8636 11178 8636 0 _095_
rlabel metal2 10166 3332 10166 3332 0 _096_
rlabel metal1 10902 8500 10902 8500 0 _097_
rlabel metal2 11362 8160 11362 8160 0 _098_
rlabel metal2 10994 7548 10994 7548 0 _099_
rlabel metal1 9706 7412 9706 7412 0 _100_
rlabel metal1 10028 8942 10028 8942 0 _101_
rlabel metal2 9338 8398 9338 8398 0 _102_
rlabel metal1 12834 3536 12834 3536 0 _103_
rlabel metal1 10580 4114 10580 4114 0 _104_
rlabel metal1 7820 8330 7820 8330 0 _105_
rlabel metal1 7038 10098 7038 10098 0 _106_
rlabel metal2 9154 11798 9154 11798 0 _107_
rlabel metal2 9246 9452 9246 9452 0 _108_
rlabel metal1 9430 7922 9430 7922 0 _109_
rlabel metal2 9522 7548 9522 7548 0 _110_
rlabel metal1 8004 6154 8004 6154 0 _111_
rlabel metal1 9108 3706 9108 3706 0 _112_
rlabel metal1 8188 3706 8188 3706 0 _113_
rlabel metal1 8004 4114 8004 4114 0 _114_
rlabel metal2 5934 4420 5934 4420 0 _115_
rlabel metal1 6302 4114 6302 4114 0 _116_
rlabel metal1 6808 3978 6808 3978 0 _117_
rlabel metal1 7406 4658 7406 4658 0 _118_
rlabel metal2 7406 4794 7406 4794 0 _119_
rlabel metal2 7498 6460 7498 6460 0 _120_
rlabel metal2 8418 11900 8418 11900 0 _121_
rlabel metal1 8556 8330 8556 8330 0 _122_
rlabel metal2 8050 6188 8050 6188 0 _123_
rlabel metal2 7406 4284 7406 4284 0 _124_
rlabel metal1 7222 4080 7222 4080 0 _125_
rlabel metal1 13754 9690 13754 9690 0 _126_
rlabel metal1 13294 11866 13294 11866 0 _127_
rlabel metal2 13662 16830 13662 16830 0 _128_
rlabel metal2 13662 14365 13662 14365 0 _129_
rlabel metal1 7820 11594 7820 11594 0 _130_
rlabel metal1 9798 8466 9798 8466 0 _131_
rlabel metal1 8878 10778 8878 10778 0 _132_
rlabel metal1 7866 11220 7866 11220 0 _133_
rlabel metal1 7682 12172 7682 12172 0 _134_
rlabel metal2 7774 11628 7774 11628 0 _135_
rlabel metal2 7590 11492 7590 11492 0 _136_
rlabel metal1 11914 11186 11914 11186 0 _137_
rlabel metal1 11638 10642 11638 10642 0 _138_
rlabel metal1 15318 11050 15318 11050 0 _139_
rlabel metal1 12236 10778 12236 10778 0 _140_
rlabel metal1 8510 11832 8510 11832 0 _141_
rlabel metal2 13202 4335 13202 4335 0 _142_
rlabel metal1 7636 11866 7636 11866 0 _143_
rlabel metal1 7176 14790 7176 14790 0 _144_
rlabel metal2 9890 16966 9890 16966 0 _145_
rlabel metal2 7222 12274 7222 12274 0 _146_
rlabel metal2 7222 11968 7222 11968 0 _147_
rlabel metal1 6992 4114 6992 4114 0 _148_
rlabel metal2 13754 8908 13754 8908 0 _149_
rlabel metal1 13570 8058 13570 8058 0 _150_
rlabel metal2 12190 6528 12190 6528 0 _151_
rlabel metal1 13110 7276 13110 7276 0 _152_
rlabel metal1 13524 7310 13524 7310 0 _153_
rlabel metal2 14122 11424 14122 11424 0 _154_
rlabel metal2 13846 11322 13846 11322 0 _155_
rlabel metal2 13110 3553 13110 3553 0 _156_
rlabel metal2 13754 12988 13754 12988 0 _157_
rlabel metal2 13938 11866 13938 11866 0 _158_
rlabel metal2 13570 9452 13570 9452 0 _159_
rlabel metal1 15502 8432 15502 8432 0 _160_
rlabel metal1 12742 14382 12742 14382 0 _161_
rlabel metal2 14858 10268 14858 10268 0 _162_
rlabel metal2 13938 7820 13938 7820 0 _163_
rlabel metal1 14399 7854 14399 7854 0 _164_
rlabel metal1 13294 7378 13294 7378 0 _165_
rlabel metal1 15134 8500 15134 8500 0 _166_
rlabel metal1 14858 8602 14858 8602 0 _167_
rlabel metal1 14306 8500 14306 8500 0 _168_
rlabel metal2 14490 8772 14490 8772 0 _169_
rlabel metal2 10902 5882 10902 5882 0 _170_
rlabel metal1 10764 5678 10764 5678 0 _171_
rlabel metal1 11454 5882 11454 5882 0 _172_
rlabel metal2 14306 10812 14306 10812 0 _173_
rlabel metal2 14122 9146 14122 9146 0 _174_
rlabel metal2 14214 8432 14214 8432 0 _175_
rlabel metal1 9706 14042 9706 14042 0 _176_
rlabel metal1 9798 14348 9798 14348 0 _177_
rlabel metal1 11592 17510 11592 17510 0 _178_
rlabel metal2 11638 15436 11638 15436 0 _179_
rlabel metal1 12880 13430 12880 13430 0 _180_
rlabel metal2 12742 14620 12742 14620 0 _181_
rlabel metal2 13018 14756 13018 14756 0 _182_
rlabel metal2 14306 15300 14306 15300 0 _183_
rlabel metal1 16698 13872 16698 13872 0 _184_
rlabel metal2 15502 12988 15502 12988 0 _185_
rlabel metal1 13524 14518 13524 14518 0 _186_
rlabel metal1 11500 14042 11500 14042 0 _187_
rlabel metal2 12558 14790 12558 14790 0 _188_
rlabel metal2 12006 16388 12006 16388 0 _189_
rlabel metal2 12190 17918 12190 17918 0 _190_
rlabel metal2 12374 18020 12374 18020 0 _191_
rlabel metal2 6486 14960 6486 14960 0 _192_
rlabel metal1 2162 14042 2162 14042 0 _193_
rlabel metal2 3266 14246 3266 14246 0 _194_
rlabel metal1 1518 13396 1518 13396 0 _195_
rlabel metal1 2530 13396 2530 13396 0 _196_
rlabel metal1 5382 6358 5382 6358 0 _197_
rlabel metal1 6532 12818 6532 12818 0 _198_
rlabel metal2 4140 12716 4140 12716 0 _199_
rlabel metal2 3358 13226 3358 13226 0 _200_
rlabel metal1 5382 5678 5382 5678 0 _201_
rlabel metal1 11178 4488 11178 4488 0 _202_
rlabel metal1 5382 5746 5382 5746 0 _203_
rlabel metal2 4830 6035 4830 6035 0 _204_
rlabel metal1 6315 12886 6315 12886 0 _205_
rlabel metal2 6394 13124 6394 13124 0 _206_
rlabel metal1 4416 13226 4416 13226 0 _207_
rlabel metal1 2392 12886 2392 12886 0 _208_
rlabel metal1 2668 12954 2668 12954 0 _209_
rlabel metal1 2208 13362 2208 13362 0 _210_
rlabel metal2 1978 13056 1978 13056 0 _211_
rlabel metal2 13570 3570 13570 3570 0 _212_
rlabel metal1 13432 3026 13432 3026 0 _213_
rlabel metal1 13156 3094 13156 3094 0 _214_
rlabel metal1 12374 5202 12374 5202 0 _215_
rlabel metal2 12006 4352 12006 4352 0 _216_
rlabel metal2 12512 4998 12512 4998 0 _217_
rlabel metal1 14030 5032 14030 5032 0 _218_
rlabel metal2 12466 9758 12466 9758 0 _219_
rlabel metal1 13294 5542 13294 5542 0 _220_
rlabel metal1 15226 5168 15226 5168 0 _221_
rlabel metal1 15456 5202 15456 5202 0 _222_
rlabel metal1 14490 5168 14490 5168 0 _223_
rlabel metal1 13925 5338 13925 5338 0 _224_
rlabel metal1 13166 3026 13166 3026 0 _225_
rlabel metal1 12834 5338 12834 5338 0 _226_
rlabel metal1 14214 5338 14214 5338 0 _227_
rlabel metal2 13110 4726 13110 4726 0 _228_
rlabel metal2 12926 4046 12926 4046 0 _229_
rlabel metal1 7728 9146 7728 9146 0 _230_
rlabel metal2 7314 9724 7314 9724 0 _231_
rlabel metal2 7084 9418 7084 9418 0 _232_
rlabel metal1 5658 10778 5658 10778 0 _233_
rlabel metal1 6992 10778 6992 10778 0 _234_
rlabel metal1 5474 11220 5474 11220 0 _235_
rlabel metal1 2346 14416 2346 14416 0 _236_
rlabel metal1 9982 12716 9982 12716 0 _237_
rlabel metal1 7912 12614 7912 12614 0 _238_
rlabel metal1 2714 12410 2714 12410 0 _239_
rlabel metal2 2438 14688 2438 14688 0 _240_
rlabel metal1 3910 11322 3910 11322 0 _241_
rlabel metal1 4370 14416 4370 14416 0 _242_
rlabel metal2 4278 15164 4278 15164 0 _243_
rlabel metal1 2346 15028 2346 15028 0 _244_
rlabel metal1 5244 14042 5244 14042 0 _245_
rlabel metal1 2622 14314 2622 14314 0 _246_
rlabel metal2 1978 14688 1978 14688 0 _247_
rlabel metal1 1978 14926 1978 14926 0 _248_
rlabel metal1 4094 8976 4094 8976 0 _249_
rlabel metal1 2530 9996 2530 9996 0 _250_
rlabel metal1 2576 10098 2576 10098 0 _251_
rlabel metal2 2530 9724 2530 9724 0 _252_
rlabel metal1 4048 10098 4048 10098 0 _253_
rlabel metal1 4462 9588 4462 9588 0 _254_
rlabel metal2 4278 9792 4278 9792 0 _255_
rlabel metal2 6486 9146 6486 9146 0 _256_
rlabel metal2 6578 9418 6578 9418 0 _257_
rlabel metal1 2898 9146 2898 9146 0 _258_
rlabel metal1 6854 10506 6854 10506 0 _259_
rlabel metal1 3174 7514 3174 7514 0 _260_
rlabel metal1 10902 3366 10902 3366 0 _261_
rlabel metal1 4830 10710 4830 10710 0 _262_
rlabel metal2 4278 10166 4278 10166 0 _263_
rlabel metal1 2898 9588 2898 9588 0 _264_
rlabel metal1 1702 9588 1702 9588 0 _265_
rlabel metal1 3036 9690 3036 9690 0 _266_
rlabel metal2 2806 9554 2806 9554 0 _267_
rlabel metal2 2346 9316 2346 9316 0 _268_
rlabel metal2 10902 3332 10902 3332 0 _269_
rlabel metal1 9522 3468 9522 3468 0 _270_
rlabel metal2 9338 3196 9338 3196 0 _271_
rlabel metal1 10166 8500 10166 8500 0 _272_
rlabel metal1 12282 10064 12282 10064 0 _273_
rlabel metal2 10258 9180 10258 9180 0 _274_
rlabel metal1 9062 6256 9062 6256 0 _275_
rlabel metal1 9568 5882 9568 5882 0 _276_
rlabel metal1 9614 6426 9614 6426 0 _277_
rlabel metal1 9246 2992 9246 2992 0 _278_
rlabel metal1 9798 3706 9798 3706 0 _279_
rlabel metal1 9476 3910 9476 3910 0 _280_
rlabel metal1 9936 2618 9936 2618 0 _281_
rlabel metal1 9982 3060 9982 3060 0 _282_
rlabel metal1 9568 4998 9568 4998 0 _283_
rlabel metal1 9016 15878 9016 15878 0 _284_
rlabel metal2 8234 5508 8234 5508 0 _285_
rlabel metal1 7866 5746 7866 5746 0 _286_
rlabel metal2 5382 6460 5382 6460 0 _287_
rlabel metal1 8142 5848 8142 5848 0 _288_
rlabel metal1 3542 5882 3542 5882 0 _289_
rlabel metal1 12880 5882 12880 5882 0 _290_
rlabel metal2 13478 9350 13478 9350 0 _291_
rlabel metal2 13018 5865 13018 5865 0 _292_
rlabel metal2 7682 6460 7682 6460 0 _293_
rlabel metal1 6394 14790 6394 14790 0 _294_
rlabel metal1 4508 6290 4508 6290 0 _295_
rlabel metal2 3818 6732 3818 6732 0 _296_
rlabel metal1 3236 6358 3236 6358 0 _297_
rlabel metal1 4048 5882 4048 5882 0 _298_
rlabel metal1 4186 6222 4186 6222 0 _299_
rlabel metal1 4048 5338 4048 5338 0 _300_
rlabel via1 3926 5678 3926 5678 0 _301_
rlabel metal1 4002 5576 4002 5576 0 _302_
rlabel metal1 10810 15096 10810 15096 0 _303_
rlabel metal1 10856 13498 10856 13498 0 _304_
rlabel metal1 10534 15028 10534 15028 0 _305_
rlabel metal1 15686 14382 15686 14382 0 _306_
rlabel metal1 15134 10778 15134 10778 0 _307_
rlabel metal2 15318 13124 15318 13124 0 _308_
rlabel metal1 16882 13838 16882 13838 0 _309_
rlabel metal1 15364 13498 15364 13498 0 _310_
rlabel metal1 14996 14382 14996 14382 0 _311_
rlabel metal1 17250 13940 17250 13940 0 _312_
rlabel metal2 17066 14144 17066 14144 0 _313_
rlabel metal2 16974 14518 16974 14518 0 _314_
rlabel metal2 15686 14620 15686 14620 0 _315_
rlabel metal1 4370 16626 4370 16626 0 _316_
rlabel metal2 5658 16456 5658 16456 0 _317_
rlabel metal1 4002 16660 4002 16660 0 _318_
rlabel metal1 6578 16558 6578 16558 0 _319_
rlabel metal1 7590 14586 7590 14586 0 _320_
rlabel metal1 7590 15130 7590 15130 0 _321_
rlabel metal2 7130 16252 7130 16252 0 _322_
rlabel metal1 7498 16626 7498 16626 0 _323_
rlabel metal1 7912 16762 7912 16762 0 _324_
rlabel metal2 10902 17680 10902 17680 0 _325_
rlabel metal1 8234 18258 8234 18258 0 _326_
rlabel metal2 10442 17442 10442 17442 0 _327_
rlabel metal2 10718 18020 10718 18020 0 _328_
rlabel metal1 11224 18258 11224 18258 0 _329_
rlabel metal2 8878 17748 8878 17748 0 _330_
rlabel metal1 5796 16558 5796 16558 0 _331_
rlabel metal1 9844 18258 9844 18258 0 _332_
rlabel metal1 9108 18258 9108 18258 0 _333_
rlabel metal1 13800 17170 13800 17170 0 _334_
rlabel metal1 13294 17748 13294 17748 0 _335_
rlabel metal1 13708 17306 13708 17306 0 _336_
rlabel metal1 11086 14382 11086 14382 0 _337_
rlabel metal1 14306 3706 14306 3706 0 _338_
rlabel metal1 16560 5338 16560 5338 0 _339_
rlabel metal2 13110 9860 13110 9860 0 _340_
rlabel metal1 2576 14994 2576 14994 0 _341_
rlabel metal1 15962 3434 15962 3434 0 _342_
rlabel metal1 8510 16218 8510 16218 0 _343_
rlabel metal1 8050 8466 8050 8466 0 _344_
rlabel via2 12650 7395 12650 7395 0 _345_
rlabel metal1 17526 6426 17526 6426 0 _346_
rlabel metal2 5750 17544 5750 17544 0 _347_
rlabel metal1 8142 11118 8142 11118 0 _348_
rlabel via2 5750 6749 5750 6749 0 _349_
rlabel metal2 6854 15572 6854 15572 0 _350_
rlabel metal2 14490 5746 14490 5746 0 _351_
rlabel metal1 12742 9928 12742 9928 0 _352_
rlabel metal1 7222 5610 7222 5610 0 _353_
rlabel metal1 4968 12138 4968 12138 0 _354_
rlabel metal1 6532 10234 6532 10234 0 _355_
rlabel metal1 4232 12138 4232 12138 0 _356_
rlabel metal1 14398 3434 14398 3434 0 _357_
rlabel metal1 13685 9962 13685 9962 0 _358_
rlabel metal2 3818 12954 3818 12954 0 _359_
rlabel metal1 14444 12818 14444 12818 0 _360_
rlabel metal2 9522 5525 9522 5525 0 _361_
rlabel metal1 8142 15504 8142 15504 0 _362_
rlabel metal1 10994 10608 10994 10608 0 _363_
rlabel metal1 11408 10098 11408 10098 0 _364_
rlabel metal1 11822 12750 11822 12750 0 _365_
rlabel metal1 9108 10030 9108 10030 0 _366_
rlabel metal1 9338 5610 9338 5610 0 _367_
rlabel metal1 15318 12852 15318 12852 0 _368_
rlabel metal1 13294 12852 13294 12852 0 _369_
rlabel metal2 13202 12410 13202 12410 0 _370_
rlabel metal2 11086 12053 11086 12053 0 _371_
rlabel metal1 15548 10030 15548 10030 0 _372_
rlabel metal1 7544 5678 7544 5678 0 _373_
rlabel metal1 8602 16116 8602 16116 0 _374_
rlabel metal1 9982 13260 9982 13260 0 _375_
rlabel metal2 15318 6817 15318 6817 0 _376_
rlabel metal1 12742 6256 12742 6256 0 _377_
rlabel metal1 11316 12410 11316 12410 0 _378_
rlabel metal1 11132 12614 11132 12614 0 _379_
rlabel metal2 15686 10030 15686 10030 0 _380_
rlabel metal2 13386 4318 13386 4318 0 _381_
rlabel metal1 11684 12410 11684 12410 0 _382_
rlabel metal1 8326 13940 8326 13940 0 _383_
rlabel metal1 4370 7412 4370 7412 0 _384_
rlabel metal1 8326 13770 8326 13770 0 _385_
rlabel metal1 8970 14416 8970 14416 0 _386_
rlabel metal1 9154 13396 9154 13396 0 _387_
rlabel metal1 2346 9554 2346 9554 0 _388_
rlabel metal1 2530 13940 2530 13940 0 _389_
rlabel metal1 17572 13906 17572 13906 0 _390_
rlabel metal1 17296 15062 17296 15062 0 clk
rlabel metal2 15226 16150 15226 16150 0 clknet_0_clk
rlabel metal1 17940 14450 17940 14450 0 clknet_1_0__leaf_clk
rlabel metal1 14444 17102 14444 17102 0 clknet_1_1__leaf_clk
rlabel metal1 16698 17646 16698 17646 0 net1
rlabel metal1 6808 3910 6808 3910 0 net10
rlabel metal1 17802 7820 17802 7820 0 net11
rlabel metal2 12374 18564 12374 18564 0 net12
rlabel metal1 1610 12954 1610 12954 0 net13
rlabel metal1 13340 2414 13340 2414 0 net14
rlabel metal2 1702 14586 1702 14586 0 net15
rlabel metal2 1702 9146 1702 9146 0 net16
rlabel metal2 9798 2686 9798 2686 0 net17
rlabel metal1 4002 13328 4002 13328 0 net18
rlabel metal1 8556 12070 8556 12070 0 net19
rlabel metal2 8510 16252 8510 16252 0 net2
rlabel metal1 8188 6222 8188 6222 0 net20
rlabel metal2 2530 13345 2530 13345 0 net21
rlabel metal1 5198 7378 5198 7378 0 net22
rlabel metal1 9246 5644 9246 5644 0 net23
rlabel metal1 14950 12682 14950 12682 0 net24
rlabel metal1 15824 6290 15824 6290 0 net25
rlabel metal1 13478 4080 13478 4080 0 net26
rlabel metal1 4738 8942 4738 8942 0 net27
rlabel metal1 6670 12308 6670 12308 0 net28
rlabel metal2 14168 13838 14168 13838 0 net29
rlabel metal1 2231 5678 2231 5678 0 net3
rlabel metal1 2162 8942 2162 8942 0 net30
rlabel metal1 2346 17646 2346 17646 0 net31
rlabel via2 14950 15453 14950 15453 0 net32
rlabel metal1 11408 18190 11408 18190 0 net33
rlabel metal2 8050 17340 8050 17340 0 net34
rlabel metal2 9706 5916 9706 5916 0 net35
rlabel metal1 7222 10234 7222 10234 0 net36
rlabel metal1 15640 7854 15640 7854 0 net37
rlabel metal1 9338 3502 9338 3502 0 net38
rlabel metal3 9108 9724 9108 9724 0 net39
rlabel metal1 17756 13906 17756 13906 0 net4
rlabel metal1 5198 13872 5198 13872 0 net40
rlabel metal2 8878 16524 8878 16524 0 net41
rlabel metal2 13110 13090 13110 13090 0 net42
rlabel metal1 9522 15504 9522 15504 0 net43
rlabel metal1 15755 16422 15755 16422 0 net44
rlabel metal1 4048 3570 4048 3570 0 net45
rlabel metal2 5566 7140 5566 7140 0 net46
rlabel metal1 7774 14382 7774 14382 0 net47
rlabel via2 5106 15997 5106 15997 0 net48
rlabel metal2 6946 14263 6946 14263 0 net49
rlabel metal2 7590 18564 7590 18564 0 net5
rlabel metal1 12834 10064 12834 10064 0 net50
rlabel viali 14673 10030 14673 10030 0 net51
rlabel metal1 13110 11696 13110 11696 0 net52
rlabel metal2 17066 10370 17066 10370 0 net53
rlabel metal1 12696 15470 12696 15470 0 net54
rlabel metal1 3634 7854 3634 7854 0 net55
rlabel metal1 9982 4046 9982 4046 0 net56
rlabel metal2 9982 15759 9982 15759 0 net57
rlabel metal2 6670 13481 6670 13481 0 net58
rlabel metal1 13754 10098 13754 10098 0 net59
rlabel metal2 11270 18564 11270 18564 0 net6
rlabel metal1 16422 12818 16422 12818 0 net60
rlabel metal1 17112 14994 17112 14994 0 net61
rlabel metal1 5842 3502 5842 3502 0 net62
rlabel metal2 2714 11390 2714 11390 0 net63
rlabel metal1 7866 9554 7866 9554 0 net64
rlabel metal2 17066 9146 17066 9146 0 net65
rlabel metal1 16928 6698 16928 6698 0 net66
rlabel metal2 5382 3332 5382 3332 0 net67
rlabel metal2 4094 11220 4094 11220 0 net68
rlabel metal2 6762 15878 6762 15878 0 net69
rlabel metal2 9154 18428 9154 18428 0 net7
rlabel metal1 9430 14994 9430 14994 0 net70
rlabel metal1 13616 10030 13616 10030 0 net71
rlabel metal1 17112 7378 17112 7378 0 net72
rlabel metal2 10074 18564 10074 18564 0 net8
rlabel metal2 9108 5780 9108 5780 0 net9
rlabel via2 17986 15011 17986 15011 0 rst
rlabel metal2 8694 19975 8694 19975 0 sine_out[0]
rlabel metal3 1096 5508 1096 5508 0 sine_out[10]
rlabel metal2 17986 14195 17986 14195 0 sine_out[11]
rlabel metal2 8050 19975 8050 19975 0 sine_out[12]
rlabel metal1 11086 18938 11086 18938 0 sine_out[13]
rlabel metal2 9982 19975 9982 19975 0 sine_out[14]
rlabel metal2 10626 19975 10626 19975 0 sine_out[15]
rlabel metal2 9062 1520 9062 1520 0 sine_out[1]
rlabel metal2 6486 1520 6486 1520 0 sine_out[2]
rlabel metal2 17986 7633 17986 7633 0 sine_out[3]
rlabel metal1 13524 18938 13524 18938 0 sine_out[4]
rlabel metal3 1096 13668 1096 13668 0 sine_out[5]
rlabel metal2 13570 1520 13570 1520 0 sine_out[6]
rlabel metal3 751 14348 751 14348 0 sine_out[7]
rlabel metal3 866 8908 866 8908 0 sine_out[8]
rlabel metal2 9706 1520 9706 1520 0 sine_out[9]
rlabel metal1 15916 13294 15916 13294 0 tcount\[0\]
rlabel metal1 17388 11730 17388 11730 0 tcount\[1\]
rlabel metal1 16836 16150 16836 16150 0 tcount\[2\]
rlabel metal1 16422 13906 16422 13906 0 tcount\[3\]
rlabel metal2 15870 16422 15870 16422 0 tcount\[4\]
rlabel metal2 16790 17680 16790 17680 0 tcount\[5\]
rlabel metal1 15916 16558 15916 16558 0 tcount\[6\]
rlabel metal1 14076 18666 14076 18666 0 tcount\[7\]
<< properties >>
string FIXED_BBOX 0 0 19560 21704
<< end >>
