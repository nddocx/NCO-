module counter_8bit (clk,
    rst,
    sine_out);
 input clk;
 input rst;
 output [15:0] sine_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire \tcount[0] ;
 wire \tcount[1] ;
 wire \tcount[2] ;
 wire \tcount[3] ;
 wire \tcount[4] ;
 wire \tcount[5] ;
 wire \tcount[6] ;
 wire \tcount[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sky130_fd_sc_hd__inv_2 _391_ (.A(net72),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _392_ (.A(\tcount[6] ),
    .Y(_331_));
 sky130_fd_sc_hd__inv_2 _393_ (.A(net34),
    .Y(_337_));
 sky130_fd_sc_hd__inv_2 _394_ (.A(net38),
    .Y(_338_));
 sky130_fd_sc_hd__inv_2 _395_ (.A(net51),
    .Y(_339_));
 sky130_fd_sc_hd__inv_2 _396_ (.A(net64),
    .Y(_340_));
 sky130_fd_sc_hd__inv_2 _397_ (.A(net31),
    .Y(_341_));
 sky130_fd_sc_hd__inv_2 _398_ (.A(net1),
    .Y(_008_));
 sky130_fd_sc_hd__nor2_1 _399_ (.A(net71),
    .B(net65),
    .Y(_342_));
 sky130_fd_sc_hd__or2_1 _400_ (.A(net69),
    .B(net64),
    .X(_343_));
 sky130_fd_sc_hd__and2_1 _401_ (.A(net72),
    .B(net65),
    .X(_344_));
 sky130_fd_sc_hd__nand2_2 _402_ (.A(net68),
    .B(net63),
    .Y(_345_));
 sky130_fd_sc_hd__xnor2_2 _403_ (.A(net71),
    .B(net65),
    .Y(_346_));
 sky130_fd_sc_hd__inv_2 _404_ (.A(net23),
    .Y(_001_));
 sky130_fd_sc_hd__nor2_4 _405_ (.A(_331_),
    .B(net34),
    .Y(_347_));
 sky130_fd_sc_hd__nand2_2 _406_ (.A(\tcount[6] ),
    .B(_337_),
    .Y(_348_));
 sky130_fd_sc_hd__nor2_2 _407_ (.A(net55),
    .B(net62),
    .Y(_349_));
 sky130_fd_sc_hd__or2_1 _408_ (.A(net58),
    .B(net64),
    .X(_350_));
 sky130_fd_sc_hd__and2b_2 _409_ (.A_N(net67),
    .B(net55),
    .X(_351_));
 sky130_fd_sc_hd__nand2b_1 _410_ (.A_N(net71),
    .B(net59),
    .Y(_352_));
 sky130_fd_sc_hd__and2b_1 _411_ (.A_N(net55),
    .B(net62),
    .X(_353_));
 sky130_fd_sc_hd__nand2b_2 _412_ (.A_N(net57),
    .B(net63),
    .Y(_354_));
 sky130_fd_sc_hd__and2_1 _413_ (.A(net70),
    .B(net56),
    .X(_355_));
 sky130_fd_sc_hd__nand2_1 _414_ (.A(net68),
    .B(net57),
    .Y(_356_));
 sky130_fd_sc_hd__nand2b_1 _415_ (.A_N(net65),
    .B(net51),
    .Y(_357_));
 sky130_fd_sc_hd__nand2b_1 _416_ (.A_N(net61),
    .B(net51),
    .Y(_358_));
 sky130_fd_sc_hd__nand2_2 _417_ (.A(net57),
    .B(net63),
    .Y(_359_));
 sky130_fd_sc_hd__xnor2_4 _418_ (.A(net57),
    .B(net63),
    .Y(_360_));
 sky130_fd_sc_hd__o21ai_4 _419_ (.A1(net68),
    .A2(net63),
    .B1(net47),
    .Y(_361_));
 sky130_fd_sc_hd__inv_2 _420_ (.A(_361_),
    .Y(_362_));
 sky130_fd_sc_hd__nor2_2 _421_ (.A(net68),
    .B(net57),
    .Y(_363_));
 sky130_fd_sc_hd__o21ai_4 _422_ (.A1(net70),
    .A2(net56),
    .B1(net49),
    .Y(_364_));
 sky130_fd_sc_hd__nor3_1 _423_ (.A(_000_),
    .B(_339_),
    .C(_360_),
    .Y(_365_));
 sky130_fd_sc_hd__nor2_1 _424_ (.A(net59),
    .B(net23),
    .Y(_366_));
 sky130_fd_sc_hd__and2b_2 _425_ (.A_N(net65),
    .B(net59),
    .X(_367_));
 sky130_fd_sc_hd__or3b_1 _426_ (.A(net72),
    .B(net66),
    .C_N(net60),
    .X(_368_));
 sky130_fd_sc_hd__o211ai_2 _427_ (.A1(net60),
    .A2(net23),
    .B1(_368_),
    .C1(net24),
    .Y(_369_));
 sky130_fd_sc_hd__nand2_1 _428_ (.A(net42),
    .B(_369_),
    .Y(_370_));
 sky130_fd_sc_hd__and2b_2 _429_ (.A_N(net55),
    .B(net70),
    .X(_371_));
 sky130_fd_sc_hd__nand2b_4 _430_ (.A_N(net61),
    .B(net71),
    .Y(_372_));
 sky130_fd_sc_hd__and2_1 _431_ (.A(net59),
    .B(net23),
    .X(_373_));
 sky130_fd_sc_hd__and2_1 _432_ (.A(net47),
    .B(net58),
    .X(_374_));
 sky130_fd_sc_hd__nand2_1 _433_ (.A(net47),
    .B(net58),
    .Y(_375_));
 sky130_fd_sc_hd__nand2_1 _434_ (.A(net48),
    .B(_354_),
    .Y(_376_));
 sky130_fd_sc_hd__a211o_1 _435_ (.A1(net59),
    .A2(net23),
    .B1(_353_),
    .C1(net24),
    .X(_377_));
 sky130_fd_sc_hd__nor2_1 _436_ (.A(_371_),
    .B(_377_),
    .Y(_378_));
 sky130_fd_sc_hd__nor3_1 _437_ (.A(net72),
    .B(net52),
    .C(net66),
    .Y(_379_));
 sky130_fd_sc_hd__nor3b_2 _438_ (.A(net51),
    .B(net65),
    .C_N(net61),
    .Y(_380_));
 sky130_fd_sc_hd__nand2_1 _439_ (.A(net24),
    .B(_367_),
    .Y(_381_));
 sky130_fd_sc_hd__or4_1 _440_ (.A(net42),
    .B(_378_),
    .C(_379_),
    .D(_380_),
    .X(_382_));
 sky130_fd_sc_hd__o21ai_1 _441_ (.A1(_365_),
    .A2(_370_),
    .B1(_382_),
    .Y(_383_));
 sky130_fd_sc_hd__and3b_1 _442_ (.A_N(net48),
    .B(net57),
    .C(net63),
    .X(_384_));
 sky130_fd_sc_hd__nor2_1 _443_ (.A(net40),
    .B(_384_),
    .Y(_385_));
 sky130_fd_sc_hd__nor2_1 _444_ (.A(net69),
    .B(net44),
    .Y(_386_));
 sky130_fd_sc_hd__o22a_1 _445_ (.A1(net22),
    .A2(_361_),
    .B1(_385_),
    .B2(_386_),
    .X(_387_));
 sky130_fd_sc_hd__nor2_4 _446_ (.A(\tcount[6] ),
    .B(net33),
    .Y(_388_));
 sky130_fd_sc_hd__or2_1 _447_ (.A(\tcount[6] ),
    .B(net33),
    .X(_389_));
 sky130_fd_sc_hd__a21bo_2 _448_ (.A1(net72),
    .A2(net66),
    .B1_N(net60),
    .X(_390_));
 sky130_fd_sc_hd__nand2_1 _449_ (.A(net24),
    .B(_390_),
    .Y(_016_));
 sky130_fd_sc_hd__a31o_1 _450_ (.A1(net42),
    .A2(_375_),
    .A3(_016_),
    .B1(net21),
    .X(_017_));
 sky130_fd_sc_hd__o21ba_2 _451_ (.A1(net55),
    .A2(net62),
    .B1_N(net45),
    .X(_018_));
 sky130_fd_sc_hd__o21bai_2 _452_ (.A1(net56),
    .A2(net62),
    .B1_N(net46),
    .Y(_019_));
 sky130_fd_sc_hd__nor2_1 _453_ (.A(net19),
    .B(_019_),
    .Y(_020_));
 sky130_fd_sc_hd__and2b_1 _454_ (.A_N(net66),
    .B(net71),
    .X(_021_));
 sky130_fd_sc_hd__nand2b_2 _455_ (.A_N(net62),
    .B(net67),
    .Y(_022_));
 sky130_fd_sc_hd__nand2_1 _456_ (.A(net52),
    .B(_355_),
    .Y(_023_));
 sky130_fd_sc_hd__nor2_1 _457_ (.A(_375_),
    .B(_022_),
    .Y(_024_));
 sky130_fd_sc_hd__nor2_1 _458_ (.A(_351_),
    .B(_371_),
    .Y(_025_));
 sky130_fd_sc_hd__xor2_4 _459_ (.A(net67),
    .B(net55),
    .X(_026_));
 sky130_fd_sc_hd__or2_1 _460_ (.A(net64),
    .B(_026_),
    .X(_027_));
 sky130_fd_sc_hd__nor2_1 _461_ (.A(net50),
    .B(_353_),
    .Y(_028_));
 sky130_fd_sc_hd__a21oi_2 _462_ (.A1(net25),
    .A2(_354_),
    .B1(net41),
    .Y(_029_));
 sky130_fd_sc_hd__nand2_1 _463_ (.A(_027_),
    .B(_029_),
    .Y(_030_));
 sky130_fd_sc_hd__nor2_4 _464_ (.A(_331_),
    .B(_337_),
    .Y(_031_));
 sky130_fd_sc_hd__nand2_4 _465_ (.A(\tcount[6] ),
    .B(net33),
    .Y(_032_));
 sky130_fd_sc_hd__o41a_1 _466_ (.A1(net27),
    .A2(_366_),
    .A3(_020_),
    .A4(_024_),
    .B1(_031_),
    .X(_033_));
 sky130_fd_sc_hd__a2bb2o_1 _467_ (.A1_N(_387_),
    .A2_N(_017_),
    .B1(_030_),
    .B2(_033_),
    .X(_034_));
 sky130_fd_sc_hd__or3_1 _468_ (.A(net69),
    .B(net57),
    .C(net64),
    .X(_035_));
 sky130_fd_sc_hd__and3b_1 _469_ (.A_N(net59),
    .B(net65),
    .C(net71),
    .X(_036_));
 sky130_fd_sc_hd__nand3b_2 _470_ (.A_N(net59),
    .B(net65),
    .C(net71),
    .Y(_037_));
 sky130_fd_sc_hd__nand2_1 _471_ (.A(_390_),
    .B(net20),
    .Y(_002_));
 sky130_fd_sc_hd__and3_1 _472_ (.A(_390_),
    .B(_035_),
    .C(_037_),
    .X(_038_));
 sky130_fd_sc_hd__nand2_1 _473_ (.A(net46),
    .B(net64),
    .Y(_039_));
 sky130_fd_sc_hd__nand2_1 _474_ (.A(_375_),
    .B(_039_),
    .Y(_040_));
 sky130_fd_sc_hd__a21bo_1 _475_ (.A1(net67),
    .A2(net62),
    .B1_N(net45),
    .X(_041_));
 sky130_fd_sc_hd__nand2_2 _476_ (.A(net51),
    .B(_372_),
    .Y(_042_));
 sky130_fd_sc_hd__a21oi_1 _477_ (.A1(net19),
    .A2(_040_),
    .B1(_038_),
    .Y(_043_));
 sky130_fd_sc_hd__and3_1 _478_ (.A(net48),
    .B(net63),
    .C(_363_),
    .X(_044_));
 sky130_fd_sc_hd__nor3b_4 _479_ (.A(net57),
    .B(net63),
    .C_N(net68),
    .Y(_045_));
 sky130_fd_sc_hd__nor2_1 _480_ (.A(net48),
    .B(_045_),
    .Y(_046_));
 sky130_fd_sc_hd__nor3_1 _481_ (.A(net45),
    .B(_351_),
    .C(_045_),
    .Y(_047_));
 sky130_fd_sc_hd__and2_1 _482_ (.A(_359_),
    .B(net18),
    .X(_048_));
 sky130_fd_sc_hd__a21o_1 _483_ (.A1(net60),
    .A2(_346_),
    .B1(_339_),
    .X(_049_));
 sky130_fd_sc_hd__or3b_1 _484_ (.A(net27),
    .B(_048_),
    .C_N(_049_),
    .X(_050_));
 sky130_fd_sc_hd__nor2_4 _485_ (.A(\tcount[6] ),
    .B(_337_),
    .Y(_051_));
 sky130_fd_sc_hd__nand2_4 _486_ (.A(_331_),
    .B(net34),
    .Y(_052_));
 sky130_fd_sc_hd__o311a_1 _487_ (.A1(net41),
    .A2(_043_),
    .A3(_044_),
    .B1(_050_),
    .C1(_051_),
    .X(_053_));
 sky130_fd_sc_hd__a211o_1 _488_ (.A1(_347_),
    .A2(_383_),
    .B1(_034_),
    .C1(_053_),
    .X(net2));
 sky130_fd_sc_hd__a221oi_1 _489_ (.A1(_000_),
    .A2(_380_),
    .B1(_038_),
    .B2(net47),
    .C1(_032_),
    .Y(_054_));
 sky130_fd_sc_hd__a32o_1 _490_ (.A1(_345_),
    .A2(_018_),
    .A3(_025_),
    .B1(_036_),
    .B2(net50),
    .X(_055_));
 sky130_fd_sc_hd__nor2_1 _491_ (.A(_342_),
    .B(_390_),
    .Y(_056_));
 sky130_fd_sc_hd__nand2_1 _492_ (.A(net56),
    .B(net19),
    .Y(_057_));
 sky130_fd_sc_hd__nor2_1 _493_ (.A(_349_),
    .B(_042_),
    .Y(_058_));
 sky130_fd_sc_hd__and2_1 _494_ (.A(net25),
    .B(net22),
    .X(_059_));
 sky130_fd_sc_hd__and3_1 _495_ (.A(_339_),
    .B(net22),
    .C(_022_),
    .X(_060_));
 sky130_fd_sc_hd__a31oi_1 _496_ (.A1(_372_),
    .A2(_040_),
    .A3(_057_),
    .B1(_060_),
    .Y(_061_));
 sky130_fd_sc_hd__a221o_1 _497_ (.A1(_347_),
    .A2(_055_),
    .B1(_061_),
    .B2(_051_),
    .C1(_054_),
    .X(_062_));
 sky130_fd_sc_hd__nand2_2 _498_ (.A(net53),
    .B(_360_),
    .Y(_063_));
 sky130_fd_sc_hd__nor2_1 _499_ (.A(net52),
    .B(net60),
    .Y(_064_));
 sky130_fd_sc_hd__or2_2 _500_ (.A(net52),
    .B(net61),
    .X(_065_));
 sky130_fd_sc_hd__nand2b_1 _501_ (.A_N(net46),
    .B(net67),
    .Y(_066_));
 sky130_fd_sc_hd__nor2_2 _502_ (.A(_345_),
    .B(_065_),
    .Y(_067_));
 sky130_fd_sc_hd__a31o_1 _503_ (.A1(net67),
    .A2(net46),
    .A3(net22),
    .B1(_067_),
    .X(_068_));
 sky130_fd_sc_hd__o21ba_1 _504_ (.A1(net56),
    .A2(net62),
    .B1_N(net67),
    .X(_069_));
 sky130_fd_sc_hd__o21bai_1 _505_ (.A1(net55),
    .A2(net62),
    .B1_N(net67),
    .Y(_070_));
 sky130_fd_sc_hd__nand2_1 _506_ (.A(net45),
    .B(_070_),
    .Y(_071_));
 sky130_fd_sc_hd__nand2_2 _507_ (.A(net62),
    .B(_026_),
    .Y(_072_));
 sky130_fd_sc_hd__a21bo_1 _508_ (.A1(net25),
    .A2(_072_),
    .B1_N(_071_),
    .X(_073_));
 sky130_fd_sc_hd__a21oi_1 _509_ (.A1(net57),
    .A2(net19),
    .B1(_364_),
    .Y(_074_));
 sky130_fd_sc_hd__a21o_1 _510_ (.A1(net56),
    .A2(net19),
    .B1(_364_),
    .X(_075_));
 sky130_fd_sc_hd__o21ba_4 _511_ (.A1(net71),
    .A2(net65),
    .B1_N(net51),
    .X(_076_));
 sky130_fd_sc_hd__nand2_1 _512_ (.A(net22),
    .B(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__a21oi_1 _513_ (.A1(_075_),
    .A2(_077_),
    .B1(_348_),
    .Y(_078_));
 sky130_fd_sc_hd__a221o_1 _514_ (.A1(_051_),
    .A2(_068_),
    .B1(_073_),
    .B2(_031_),
    .C1(net26),
    .X(_079_));
 sky130_fd_sc_hd__o22a_1 _515_ (.A1(net36),
    .A2(_062_),
    .B1(_078_),
    .B2(_079_),
    .X(_080_));
 sky130_fd_sc_hd__a21o_1 _516_ (.A1(net65),
    .A2(_351_),
    .B1(_364_),
    .X(_081_));
 sky130_fd_sc_hd__and3b_1 _517_ (.A_N(net53),
    .B(net60),
    .C(net72),
    .X(_082_));
 sky130_fd_sc_hd__nor2_1 _518_ (.A(net37),
    .B(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__o211a_1 _519_ (.A1(net51),
    .A2(_021_),
    .B1(_376_),
    .C1(net37),
    .X(_084_));
 sky130_fd_sc_hd__a211oi_1 _520_ (.A1(_081_),
    .A2(_083_),
    .B1(_084_),
    .C1(net21),
    .Y(_085_));
 sky130_fd_sc_hd__or3_1 _521_ (.A(net51),
    .B(_360_),
    .C(_021_),
    .X(_086_));
 sky130_fd_sc_hd__nor2_1 _522_ (.A(_349_),
    .B(_364_),
    .Y(_087_));
 sky130_fd_sc_hd__o311a_1 _523_ (.A1(_349_),
    .A2(_355_),
    .A3(_364_),
    .B1(_086_),
    .C1(net29),
    .X(_088_));
 sky130_fd_sc_hd__and3_1 _524_ (.A(net69),
    .B(net58),
    .C(net63),
    .X(_089_));
 sky130_fd_sc_hd__nor2_1 _525_ (.A(net47),
    .B(_089_),
    .Y(_090_));
 sky130_fd_sc_hd__a31o_1 _526_ (.A1(net68),
    .A2(net57),
    .A3(net63),
    .B1(net48),
    .X(_091_));
 sky130_fd_sc_hd__or2_1 _527_ (.A(_045_),
    .B(_091_),
    .X(_092_));
 sky130_fd_sc_hd__o31a_1 _528_ (.A1(net24),
    .A2(_351_),
    .A3(_021_),
    .B1(net38),
    .X(_093_));
 sky130_fd_sc_hd__o21a_1 _529_ (.A1(_069_),
    .A2(_092_),
    .B1(_093_),
    .X(_094_));
 sky130_fd_sc_hd__a311o_1 _530_ (.A1(net50),
    .A2(_340_),
    .A3(_363_),
    .B1(_380_),
    .C1(_344_),
    .X(_095_));
 sky130_fd_sc_hd__nor2_1 _531_ (.A(_357_),
    .B(_371_),
    .Y(_096_));
 sky130_fd_sc_hd__o211a_1 _532_ (.A1(_344_),
    .A2(_026_),
    .B1(_039_),
    .C1(net37),
    .X(_097_));
 sky130_fd_sc_hd__a211o_1 _533_ (.A1(net29),
    .A2(_095_),
    .B1(_097_),
    .C1(_052_),
    .X(_098_));
 sky130_fd_sc_hd__o311a_1 _534_ (.A1(_032_),
    .A2(_088_),
    .A3(_094_),
    .B1(_098_),
    .C1(net30),
    .X(_099_));
 sky130_fd_sc_hd__inv_2 _535_ (.A(_099_),
    .Y(_100_));
 sky130_fd_sc_hd__and3_1 _536_ (.A(net47),
    .B(_027_),
    .C(_072_),
    .X(_101_));
 sky130_fd_sc_hd__a211o_1 _537_ (.A1(net71),
    .A2(_380_),
    .B1(_101_),
    .C1(net37),
    .X(_102_));
 sky130_fd_sc_hd__a21o_1 _538_ (.A1(net50),
    .A2(_349_),
    .B1(net26),
    .X(_103_));
 sky130_fd_sc_hd__a21o_1 _539_ (.A1(_026_),
    .A2(_028_),
    .B1(_103_),
    .X(_104_));
 sky130_fd_sc_hd__nand2_1 _540_ (.A(_385_),
    .B(_066_),
    .Y(_105_));
 sky130_fd_sc_hd__a21o_1 _541_ (.A1(_000_),
    .A2(net66),
    .B1(net28),
    .X(_106_));
 sky130_fd_sc_hd__nand2_1 _542_ (.A(_375_),
    .B(_065_),
    .Y(_107_));
 sky130_fd_sc_hd__a31o_1 _543_ (.A1(_375_),
    .A2(_022_),
    .A3(_065_),
    .B1(_106_),
    .X(_108_));
 sky130_fd_sc_hd__o211a_1 _544_ (.A1(_101_),
    .A2(_105_),
    .B1(_108_),
    .C1(_347_),
    .X(_109_));
 sky130_fd_sc_hd__a31o_1 _545_ (.A1(_388_),
    .A2(_102_),
    .A3(_104_),
    .B1(_109_),
    .X(_110_));
 sky130_fd_sc_hd__o32a_1 _546_ (.A1(net30),
    .A2(_080_),
    .A3(_085_),
    .B1(_100_),
    .B2(_110_),
    .X(net9));
 sky130_fd_sc_hd__nand2_1 _547_ (.A(net22),
    .B(_372_),
    .Y(_111_));
 sky130_fd_sc_hd__a21oi_1 _548_ (.A1(net20),
    .A2(_111_),
    .B1(net46),
    .Y(_112_));
 sky130_fd_sc_hd__o21ai_1 _549_ (.A1(_096_),
    .A2(_112_),
    .B1(net35),
    .Y(_113_));
 sky130_fd_sc_hd__a21o_1 _550_ (.A1(net46),
    .A2(_111_),
    .B1(_105_),
    .X(_114_));
 sky130_fd_sc_hd__or3_1 _551_ (.A(net45),
    .B(net19),
    .C(_353_),
    .X(_115_));
 sky130_fd_sc_hd__or2_1 _552_ (.A(_351_),
    .B(_041_),
    .X(_116_));
 sky130_fd_sc_hd__a21oi_1 _553_ (.A1(_115_),
    .A2(_116_),
    .B1(net35),
    .Y(_117_));
 sky130_fd_sc_hd__a41o_1 _554_ (.A1(net35),
    .A2(_019_),
    .A3(_041_),
    .A4(_066_),
    .B1(_117_),
    .X(_118_));
 sky130_fd_sc_hd__o211a_1 _555_ (.A1(net46),
    .A2(_373_),
    .B1(_063_),
    .C1(net35),
    .X(_119_));
 sky130_fd_sc_hd__a31o_1 _556_ (.A1(_385_),
    .A2(_039_),
    .A3(_042_),
    .B1(_348_),
    .X(_120_));
 sky130_fd_sc_hd__a221o_1 _557_ (.A1(_362_),
    .A2(_390_),
    .B1(_090_),
    .B2(_343_),
    .C1(net44),
    .X(_121_));
 sky130_fd_sc_hd__nand2_1 _558_ (.A(net36),
    .B(_361_),
    .Y(_122_));
 sky130_fd_sc_hd__o311a_1 _559_ (.A1(_344_),
    .A2(_363_),
    .A3(_122_),
    .B1(_121_),
    .C1(_031_),
    .X(_123_));
 sky130_fd_sc_hd__o221ai_1 _560_ (.A1(_052_),
    .A2(_118_),
    .B1(_119_),
    .B2(_120_),
    .C1(net30),
    .Y(_124_));
 sky130_fd_sc_hd__a31o_1 _561_ (.A1(_388_),
    .A2(_113_),
    .A3(_114_),
    .B1(_123_),
    .X(_125_));
 sky130_fd_sc_hd__a21oi_1 _562_ (.A1(_357_),
    .A2(_358_),
    .B1(_045_),
    .Y(_126_));
 sky130_fd_sc_hd__nor2_1 _563_ (.A(net52),
    .B(_072_),
    .Y(_127_));
 sky130_fd_sc_hd__and4_1 _564_ (.A(net72),
    .B(net52),
    .C(net60),
    .D(\tcount[1] ),
    .X(_128_));
 sky130_fd_sc_hd__or2_1 _565_ (.A(net43),
    .B(_128_),
    .X(_129_));
 sky130_fd_sc_hd__o221a_1 _566_ (.A1(_370_),
    .A2(_126_),
    .B1(_127_),
    .B2(_129_),
    .C1(_388_),
    .X(_130_));
 sky130_fd_sc_hd__a21oi_1 _567_ (.A1(_040_),
    .A2(_057_),
    .B1(net37),
    .Y(_131_));
 sky130_fd_sc_hd__a221o_1 _568_ (.A1(_022_),
    .A2(_028_),
    .B1(_040_),
    .B2(_057_),
    .C1(net42),
    .X(_132_));
 sky130_fd_sc_hd__or3_1 _569_ (.A(net47),
    .B(_045_),
    .C(_106_),
    .X(_133_));
 sky130_fd_sc_hd__and3_1 _570_ (.A(net48),
    .B(_356_),
    .C(_359_),
    .X(_134_));
 sky130_fd_sc_hd__or3b_1 _571_ (.A(net27),
    .B(_349_),
    .C_N(_134_),
    .X(_135_));
 sky130_fd_sc_hd__a31o_1 _572_ (.A1(_132_),
    .A2(_133_),
    .A3(_135_),
    .B1(_348_),
    .X(_136_));
 sky130_fd_sc_hd__a221o_1 _573_ (.A1(net23),
    .A2(_028_),
    .B1(net20),
    .B2(net52),
    .C1(net42),
    .X(_137_));
 sky130_fd_sc_hd__or3_1 _574_ (.A(net52),
    .B(net66),
    .C(_363_),
    .X(_138_));
 sky130_fd_sc_hd__and4b_1 _575_ (.A_N(net72),
    .B(net53),
    .C(net61),
    .D(net66),
    .X(_139_));
 sky130_fd_sc_hd__or3b_1 _576_ (.A(_139_),
    .B(net28),
    .C_N(_138_),
    .X(_140_));
 sky130_fd_sc_hd__a31o_1 _577_ (.A1(_031_),
    .A2(_137_),
    .A3(_140_),
    .B1(net31),
    .X(_141_));
 sky130_fd_sc_hd__or2_2 _578_ (.A(net55),
    .B(_041_),
    .X(_142_));
 sky130_fd_sc_hd__a211o_1 _579_ (.A1(_026_),
    .A2(_040_),
    .B1(_076_),
    .C1(net41),
    .X(_143_));
 sky130_fd_sc_hd__a311o_1 _580_ (.A1(_343_),
    .A2(_350_),
    .A3(_359_),
    .B1(net47),
    .C1(net27),
    .X(_144_));
 sky130_fd_sc_hd__nand2_1 _581_ (.A(net43),
    .B(net47),
    .Y(_145_));
 sky130_fd_sc_hd__or3_1 _582_ (.A(net28),
    .B(net19),
    .C(_364_),
    .X(_146_));
 sky130_fd_sc_hd__a31o_1 _583_ (.A1(_143_),
    .A2(_144_),
    .A3(_146_),
    .B1(_052_),
    .X(_147_));
 sky130_fd_sc_hd__and4bb_1 _584_ (.A_N(_130_),
    .B_N(_141_),
    .C(_147_),
    .D(_136_),
    .X(_148_));
 sky130_fd_sc_hd__o21ba_1 _585_ (.A1(_124_),
    .A2(_125_),
    .B1_N(_148_),
    .X(net10));
 sky130_fd_sc_hd__a211o_1 _586_ (.A1(net59),
    .A2(_076_),
    .B1(_126_),
    .C1(_067_),
    .X(_149_));
 sky130_fd_sc_hd__o31a_1 _587_ (.A1(net37),
    .A2(_363_),
    .A3(_367_),
    .B1(_149_),
    .X(_150_));
 sky130_fd_sc_hd__o211a_1 _588_ (.A1(_364_),
    .A2(_373_),
    .B1(_092_),
    .C1(net38),
    .X(_151_));
 sky130_fd_sc_hd__nand2_1 _589_ (.A(_345_),
    .B(_028_),
    .Y(_152_));
 sky130_fd_sc_hd__a31o_1 _590_ (.A1(net29),
    .A2(net20),
    .A3(_152_),
    .B1(_348_),
    .X(_153_));
 sky130_fd_sc_hd__a32o_1 _591_ (.A1(net53),
    .A2(net66),
    .A3(_026_),
    .B1(_076_),
    .B2(net22),
    .X(_154_));
 sky130_fd_sc_hd__nand2_1 _592_ (.A(net43),
    .B(_154_),
    .Y(_155_));
 sky130_fd_sc_hd__a21oi_2 _593_ (.A1(net71),
    .A2(net59),
    .B1(net51),
    .Y(_156_));
 sky130_fd_sc_hd__nand2_1 _594_ (.A(net23),
    .B(_156_),
    .Y(_157_));
 sky130_fd_sc_hd__a31o_1 _595_ (.A1(_023_),
    .A2(_063_),
    .A3(_157_),
    .B1(net42),
    .X(_158_));
 sky130_fd_sc_hd__a21o_1 _596_ (.A1(_155_),
    .A2(_158_),
    .B1(net21),
    .X(_159_));
 sky130_fd_sc_hd__o31a_1 _597_ (.A1(net24),
    .A2(_045_),
    .A3(_056_),
    .B1(_083_),
    .X(_160_));
 sky130_fd_sc_hd__a21oi_1 _598_ (.A1(_368_),
    .A2(net20),
    .B1(net25),
    .Y(_161_));
 sky130_fd_sc_hd__a211o_1 _599_ (.A1(net61),
    .A2(_076_),
    .B1(_161_),
    .C1(_067_),
    .X(_162_));
 sky130_fd_sc_hd__a21oi_1 _600_ (.A1(net37),
    .A2(_162_),
    .B1(_160_),
    .Y(_163_));
 sky130_fd_sc_hd__o21a_1 _601_ (.A1(_052_),
    .A2(_150_),
    .B1(_159_),
    .X(_164_));
 sky130_fd_sc_hd__o221a_1 _602_ (.A1(_151_),
    .A2(_153_),
    .B1(_163_),
    .B2(_032_),
    .C1(net30),
    .X(_165_));
 sky130_fd_sc_hd__or2_1 _603_ (.A(_344_),
    .B(_082_),
    .X(_166_));
 sky130_fd_sc_hd__a311o_1 _604_ (.A1(net39),
    .A2(_042_),
    .A3(_166_),
    .B1(_160_),
    .C1(_032_),
    .X(_167_));
 sky130_fd_sc_hd__or2_1 _605_ (.A(net37),
    .B(_072_),
    .X(_168_));
 sky130_fd_sc_hd__a31o_1 _606_ (.A1(_051_),
    .A2(_149_),
    .A3(_168_),
    .B1(net30),
    .X(_169_));
 sky130_fd_sc_hd__o31a_1 _607_ (.A1(net24),
    .A2(_367_),
    .A3(_025_),
    .B1(_092_),
    .X(_170_));
 sky130_fd_sc_hd__a221o_1 _608_ (.A1(net50),
    .A2(net20),
    .B1(_057_),
    .B2(_372_),
    .C1(net38),
    .X(_171_));
 sky130_fd_sc_hd__o211a_1 _609_ (.A1(net29),
    .A2(_170_),
    .B1(_171_),
    .C1(_347_),
    .X(_172_));
 sky130_fd_sc_hd__o21a_1 _610_ (.A1(_000_),
    .A2(_376_),
    .B1(_065_),
    .X(_173_));
 sky130_fd_sc_hd__o211a_1 _611_ (.A1(net42),
    .A2(_173_),
    .B1(_155_),
    .C1(_388_),
    .X(_174_));
 sky130_fd_sc_hd__or3b_1 _612_ (.A(_169_),
    .B(_172_),
    .C_N(_167_),
    .X(_175_));
 sky130_fd_sc_hd__o2bb2a_1 _613_ (.A1_N(_164_),
    .A2_N(_165_),
    .B1(_174_),
    .B2(_175_),
    .X(net11));
 sky130_fd_sc_hd__nor2_1 _614_ (.A(_027_),
    .B(_107_),
    .Y(_176_));
 sky130_fd_sc_hd__or3b_1 _615_ (.A(net25),
    .B(net22),
    .C_N(_386_),
    .X(_177_));
 sky130_fd_sc_hd__o211a_1 _616_ (.A1(net28),
    .A2(_176_),
    .B1(_177_),
    .C1(_388_),
    .X(_178_));
 sky130_fd_sc_hd__nand2_1 _617_ (.A(_345_),
    .B(_064_),
    .Y(_179_));
 sky130_fd_sc_hd__o21a_1 _618_ (.A1(net60),
    .A2(net23),
    .B1(_156_),
    .X(_180_));
 sky130_fd_sc_hd__a31o_1 _619_ (.A1(net72),
    .A2(net52),
    .A3(net60),
    .B1(net43),
    .X(_181_));
 sky130_fd_sc_hd__o32ai_1 _620_ (.A1(net28),
    .A2(_060_),
    .A3(_161_),
    .B1(_180_),
    .B2(_181_),
    .Y(_182_));
 sky130_fd_sc_hd__nor2_1 _621_ (.A(_379_),
    .B(_064_),
    .Y(_183_));
 sky130_fd_sc_hd__a31o_1 _622_ (.A1(net29),
    .A2(_377_),
    .A3(_183_),
    .B1(net33),
    .X(_184_));
 sky130_fd_sc_hd__nor4_1 _623_ (.A(net28),
    .B(_380_),
    .C(_082_),
    .D(_139_),
    .Y(_185_));
 sky130_fd_sc_hd__a311o_1 _624_ (.A1(net29),
    .A2(_377_),
    .A3(_183_),
    .B1(_185_),
    .C1(net33),
    .X(_186_));
 sky130_fd_sc_hd__a21bo_1 _625_ (.A1(net60),
    .A2(_076_),
    .B1_N(_364_),
    .X(_187_));
 sky130_fd_sc_hd__a221o_1 _626_ (.A1(_029_),
    .A2(_049_),
    .B1(_187_),
    .B2(net43),
    .C1(_337_),
    .X(_188_));
 sky130_fd_sc_hd__a32o_1 _627_ (.A1(\tcount[6] ),
    .A2(_186_),
    .A3(_188_),
    .B1(_051_),
    .B2(_182_),
    .X(_189_));
 sky130_fd_sc_hd__a21oi_1 _628_ (.A1(_178_),
    .A2(_179_),
    .B1(_189_),
    .Y(_190_));
 sky130_fd_sc_hd__or3_1 _629_ (.A(net31),
    .B(_178_),
    .C(_189_),
    .X(_191_));
 sky130_fd_sc_hd__o21ai_1 _630_ (.A1(_341_),
    .A2(_190_),
    .B1(_191_),
    .Y(net12));
 sky130_fd_sc_hd__o22a_1 _631_ (.A1(net69),
    .A2(net22),
    .B1(_361_),
    .B2(_089_),
    .X(_192_));
 sky130_fd_sc_hd__o21ai_1 _632_ (.A1(_044_),
    .A2(_192_),
    .B1(net40),
    .Y(_193_));
 sky130_fd_sc_hd__a31o_1 _633_ (.A1(net47),
    .A2(_343_),
    .A3(_037_),
    .B1(net40),
    .X(_194_));
 sky130_fd_sc_hd__or2_1 _634_ (.A(net18),
    .B(_194_),
    .X(_195_));
 sky130_fd_sc_hd__a21oi_1 _635_ (.A1(_193_),
    .A2(_195_),
    .B1(net21),
    .Y(_196_));
 sky130_fd_sc_hd__o211a_1 _636_ (.A1(net68),
    .A2(net22),
    .B1(_022_),
    .C1(_356_),
    .X(_197_));
 sky130_fd_sc_hd__a221o_1 _637_ (.A1(net68),
    .A2(_354_),
    .B1(_359_),
    .B2(_069_),
    .C1(net48),
    .X(_198_));
 sky130_fd_sc_hd__a311o_1 _638_ (.A1(_354_),
    .A2(_356_),
    .A3(_198_),
    .B1(_067_),
    .C1(net28),
    .X(_199_));
 sky130_fd_sc_hd__o311a_1 _639_ (.A1(net41),
    .A2(_048_),
    .A3(_058_),
    .B1(_199_),
    .C1(_031_),
    .X(_200_));
 sky130_fd_sc_hd__o311a_1 _640_ (.A1(net45),
    .A2(_353_),
    .A3(_025_),
    .B1(_361_),
    .C1(net35),
    .X(_201_));
 sky130_fd_sc_hd__or3_1 _641_ (.A(net24),
    .B(_351_),
    .C(_036_),
    .X(_202_));
 sky130_fd_sc_hd__a21oi_1 _642_ (.A1(_115_),
    .A2(_202_),
    .B1(net35),
    .Y(_203_));
 sky130_fd_sc_hd__o21a_1 _643_ (.A1(_201_),
    .A2(_203_),
    .B1(_347_),
    .X(_204_));
 sky130_fd_sc_hd__o21a_1 _644_ (.A1(_355_),
    .A2(_361_),
    .B1(net28),
    .X(_205_));
 sky130_fd_sc_hd__a32o_1 _645_ (.A1(net41),
    .A2(_063_),
    .A3(_198_),
    .B1(_205_),
    .B2(_369_),
    .X(_206_));
 sky130_fd_sc_hd__nand2_1 _646_ (.A(_051_),
    .B(_206_),
    .Y(_207_));
 sky130_fd_sc_hd__or4b_1 _647_ (.A(_196_),
    .B(_200_),
    .C(_204_),
    .D_N(_207_),
    .X(_208_));
 sky130_fd_sc_hd__a21o_1 _648_ (.A1(net68),
    .A2(_018_),
    .B1(_194_),
    .X(_209_));
 sky130_fd_sc_hd__a21o_1 _649_ (.A1(_193_),
    .A2(_209_),
    .B1(_389_),
    .X(_210_));
 sky130_fd_sc_hd__and4bb_1 _650_ (.A_N(_200_),
    .B_N(_204_),
    .C(_207_),
    .D(_210_),
    .X(_211_));
 sky130_fd_sc_hd__mux2_1 _651_ (.A0(_208_),
    .A1(_211_),
    .S(_341_),
    .X(net13));
 sky130_fd_sc_hd__a21oi_1 _652_ (.A1(net66),
    .A2(_156_),
    .B1(_103_),
    .Y(_212_));
 sky130_fd_sc_hd__o21a_1 _653_ (.A1(_087_),
    .A2(_112_),
    .B1(net26),
    .X(_213_));
 sky130_fd_sc_hd__o21ai_1 _654_ (.A1(_212_),
    .A2(_213_),
    .B1(_388_),
    .Y(_214_));
 sky130_fd_sc_hd__o211a_1 _655_ (.A1(net50),
    .A2(_366_),
    .B1(_377_),
    .C1(net38),
    .X(_215_));
 sky130_fd_sc_hd__nand2_1 _656_ (.A(net20),
    .B(_076_),
    .Y(_216_));
 sky130_fd_sc_hd__and3_1 _657_ (.A(net26),
    .B(_202_),
    .C(_216_),
    .X(_217_));
 sky130_fd_sc_hd__or3_1 _658_ (.A(_032_),
    .B(_215_),
    .C(_217_),
    .X(_218_));
 sky130_fd_sc_hd__a32o_1 _659_ (.A1(net50),
    .A2(_352_),
    .A3(_022_),
    .B1(_358_),
    .B2(_340_),
    .X(_219_));
 sky130_fd_sc_hd__a22o_1 _660_ (.A1(_029_),
    .A2(_042_),
    .B1(_219_),
    .B2(net37),
    .X(_220_));
 sky130_fd_sc_hd__a211o_1 _661_ (.A1(net59),
    .A2(_001_),
    .B1(_036_),
    .C1(net24),
    .X(_221_));
 sky130_fd_sc_hd__a22o_1 _662_ (.A1(net51),
    .A2(_372_),
    .B1(net20),
    .B2(_076_),
    .X(_222_));
 sky130_fd_sc_hd__a22o_1 _663_ (.A1(_083_),
    .A2(_221_),
    .B1(_222_),
    .B2(net38),
    .X(_223_));
 sky130_fd_sc_hd__o2bb2a_1 _664_ (.A1_N(_051_),
    .A2_N(_220_),
    .B1(_223_),
    .B2(_348_),
    .X(_224_));
 sky130_fd_sc_hd__and3_1 _665_ (.A(net30),
    .B(_218_),
    .C(_224_),
    .X(_225_));
 sky130_fd_sc_hd__o21ai_1 _666_ (.A1(_215_),
    .A2(_217_),
    .B1(_031_),
    .Y(_226_));
 sky130_fd_sc_hd__nand2_1 _667_ (.A(_347_),
    .B(_223_),
    .Y(_227_));
 sky130_fd_sc_hd__a311o_1 _668_ (.A1(net26),
    .A2(_381_),
    .A3(_142_),
    .B1(_212_),
    .C1(net21),
    .X(_228_));
 sky130_fd_sc_hd__o2111a_1 _669_ (.A1(_052_),
    .A2(_220_),
    .B1(_226_),
    .C1(_227_),
    .D1(_228_),
    .X(_229_));
 sky130_fd_sc_hd__a22oi_1 _670_ (.A1(_214_),
    .A2(_225_),
    .B1(_229_),
    .B2(_341_),
    .Y(net14));
 sky130_fd_sc_hd__or2_1 _671_ (.A(_344_),
    .B(_364_),
    .X(_230_));
 sky130_fd_sc_hd__nand2_1 _672_ (.A(net36),
    .B(_066_),
    .Y(_231_));
 sky130_fd_sc_hd__a2bb2o_1 _673_ (.A1_N(_366_),
    .A2_N(_231_),
    .B1(_230_),
    .B2(_385_),
    .X(_232_));
 sky130_fd_sc_hd__a221o_1 _674_ (.A1(net25),
    .A2(_072_),
    .B1(_074_),
    .B2(_354_),
    .C1(net41),
    .X(_233_));
 sky130_fd_sc_hd__nor2_1 _675_ (.A(net58),
    .B(_039_),
    .Y(_234_));
 sky130_fd_sc_hd__a211o_1 _676_ (.A1(_345_),
    .A2(_107_),
    .B1(_234_),
    .C1(net27),
    .X(_235_));
 sky130_fd_sc_hd__a32o_1 _677_ (.A1(_031_),
    .A2(_233_),
    .A3(_235_),
    .B1(_232_),
    .B2(_347_),
    .X(_236_));
 sky130_fd_sc_hd__or3_1 _678_ (.A(net29),
    .B(_379_),
    .C(_380_),
    .X(_237_));
 sky130_fd_sc_hd__a31o_1 _679_ (.A1(net52),
    .A2(_027_),
    .A3(_072_),
    .B1(_237_),
    .X(_238_));
 sky130_fd_sc_hd__a311o_1 _680_ (.A1(net48),
    .A2(_354_),
    .A3(_356_),
    .B1(_046_),
    .C1(net41),
    .X(_239_));
 sky130_fd_sc_hd__a31o_1 _681_ (.A1(_331_),
    .A2(_238_),
    .A3(_239_),
    .B1(_388_),
    .X(_240_));
 sky130_fd_sc_hd__o21a_1 _682_ (.A1(_045_),
    .A2(_069_),
    .B1(net48),
    .X(_241_));
 sky130_fd_sc_hd__o21ai_1 _683_ (.A1(_059_),
    .A2(_241_),
    .B1(net40),
    .Y(_242_));
 sky130_fd_sc_hd__or4_1 _684_ (.A(net40),
    .B(_349_),
    .C(_363_),
    .D(_384_),
    .X(_243_));
 sky130_fd_sc_hd__a21o_1 _685_ (.A1(_242_),
    .A2(_243_),
    .B1(net34),
    .X(_244_));
 sky130_fd_sc_hd__nand2_1 _686_ (.A(_385_),
    .B(_142_),
    .Y(_245_));
 sky130_fd_sc_hd__a21o_1 _687_ (.A1(_242_),
    .A2(_245_),
    .B1(net34),
    .X(_246_));
 sky130_fd_sc_hd__a21oi_1 _688_ (.A1(_240_),
    .A2(_246_),
    .B1(_236_),
    .Y(_247_));
 sky130_fd_sc_hd__a211o_1 _689_ (.A1(_240_),
    .A2(_244_),
    .B1(_341_),
    .C1(_236_),
    .X(_248_));
 sky130_fd_sc_hd__o21ai_1 _690_ (.A1(net31),
    .A2(_247_),
    .B1(_248_),
    .Y(net15));
 sky130_fd_sc_hd__or3_1 _691_ (.A(net26),
    .B(net45),
    .C(_070_),
    .X(_249_));
 sky130_fd_sc_hd__o41a_1 _692_ (.A1(net27),
    .A2(net62),
    .A3(_363_),
    .A4(_018_),
    .B1(_249_),
    .X(_250_));
 sky130_fd_sc_hd__and3_1 _693_ (.A(net45),
    .B(_345_),
    .C(_026_),
    .X(_251_));
 sky130_fd_sc_hd__o31ai_1 _694_ (.A1(net36),
    .A2(_047_),
    .A3(_251_),
    .B1(_250_),
    .Y(_252_));
 sky130_fd_sc_hd__or3_1 _695_ (.A(net27),
    .B(net18),
    .C(_241_),
    .X(_253_));
 sky130_fd_sc_hd__a21o_1 _696_ (.A1(net25),
    .A2(_390_),
    .B1(net36),
    .X(_254_));
 sky130_fd_sc_hd__a21o_1 _697_ (.A1(net45),
    .A2(_197_),
    .B1(_254_),
    .X(_255_));
 sky130_fd_sc_hd__a31o_1 _698_ (.A1(_340_),
    .A2(_066_),
    .A3(_107_),
    .B1(net36),
    .X(_256_));
 sky130_fd_sc_hd__or3_1 _699_ (.A(net25),
    .B(_355_),
    .C(_106_),
    .X(_257_));
 sky130_fd_sc_hd__a31oi_1 _700_ (.A1(_249_),
    .A2(_256_),
    .A3(_257_),
    .B1(_052_),
    .Y(_258_));
 sky130_fd_sc_hd__a21oi_1 _701_ (.A1(_346_),
    .A2(_065_),
    .B1(_371_),
    .Y(_259_));
 sky130_fd_sc_hd__and3b_1 _702_ (.A_N(net55),
    .B(net46),
    .C(net67),
    .X(_260_));
 sky130_fd_sc_hd__o21ai_1 _703_ (.A1(_342_),
    .A2(_026_),
    .B1(net50),
    .Y(_261_));
 sky130_fd_sc_hd__a311o_1 _704_ (.A1(net48),
    .A2(_354_),
    .A3(_356_),
    .B1(_260_),
    .C1(net41),
    .X(_262_));
 sky130_fd_sc_hd__o311a_1 _705_ (.A1(net27),
    .A2(_074_),
    .A3(_259_),
    .B1(_262_),
    .C1(_347_),
    .X(_263_));
 sky130_fd_sc_hd__a31o_1 _706_ (.A1(_031_),
    .A2(_253_),
    .A3(_255_),
    .B1(_263_),
    .X(_264_));
 sky130_fd_sc_hd__a211o_1 _707_ (.A1(_388_),
    .A2(_252_),
    .B1(_258_),
    .C1(_264_),
    .X(_265_));
 sky130_fd_sc_hd__a211o_1 _708_ (.A1(net67),
    .A2(_018_),
    .B1(_251_),
    .C1(net36),
    .X(_266_));
 sky130_fd_sc_hd__a21oi_1 _709_ (.A1(_250_),
    .A2(_266_),
    .B1(net21),
    .Y(_267_));
 sky130_fd_sc_hd__or4_1 _710_ (.A(net30),
    .B(_258_),
    .C(_264_),
    .D(_267_),
    .X(_268_));
 sky130_fd_sc_hd__a21bo_1 _711_ (.A1(net30),
    .A2(_265_),
    .B1_N(_268_),
    .X(net16));
 sky130_fd_sc_hd__nand2_1 _712_ (.A(net19),
    .B(_018_),
    .Y(_269_));
 sky130_fd_sc_hd__a21o_1 _713_ (.A1(_261_),
    .A2(_269_),
    .B1(net26),
    .X(_270_));
 sky130_fd_sc_hd__o31a_1 _714_ (.A1(net38),
    .A2(_020_),
    .A3(_096_),
    .B1(_270_),
    .X(_271_));
 sky130_fd_sc_hd__a31o_1 _715_ (.A1(net36),
    .A2(_071_),
    .A3(_198_),
    .B1(_348_),
    .X(_272_));
 sky130_fd_sc_hd__o221a_1 _716_ (.A1(_355_),
    .A2(_364_),
    .B1(_069_),
    .B2(net50),
    .C1(net28),
    .X(_273_));
 sky130_fd_sc_hd__a311o_1 _717_ (.A1(net37),
    .A2(_138_),
    .A3(_142_),
    .B1(_273_),
    .C1(_052_),
    .X(_274_));
 sky130_fd_sc_hd__nand2_1 _718_ (.A(net46),
    .B(net23),
    .Y(_275_));
 sky130_fd_sc_hd__o221a_1 _719_ (.A1(_361_),
    .A2(_367_),
    .B1(_019_),
    .B2(net23),
    .C1(net35),
    .X(_276_));
 sky130_fd_sc_hd__a311o_1 _720_ (.A1(net26),
    .A2(_025_),
    .A3(_275_),
    .B1(_276_),
    .C1(_032_),
    .X(_277_));
 sky130_fd_sc_hd__o211a_1 _721_ (.A1(_131_),
    .A2(_272_),
    .B1(_274_),
    .C1(_277_),
    .X(_278_));
 sky130_fd_sc_hd__a211o_1 _722_ (.A1(_018_),
    .A2(_057_),
    .B1(_096_),
    .C1(net38),
    .X(_279_));
 sky130_fd_sc_hd__a21o_1 _723_ (.A1(_270_),
    .A2(_279_),
    .B1(net21),
    .X(_280_));
 sky130_fd_sc_hd__nand2_1 _724_ (.A(_278_),
    .B(_280_),
    .Y(_281_));
 sky130_fd_sc_hd__o211a_1 _725_ (.A1(net21),
    .A2(_271_),
    .B1(_278_),
    .C1(_341_),
    .X(_282_));
 sky130_fd_sc_hd__a21o_1 _726_ (.A1(net32),
    .A2(_281_),
    .B1(_282_),
    .X(net17));
 sky130_fd_sc_hd__o41a_1 _727_ (.A1(net50),
    .A2(_342_),
    .A3(_351_),
    .A4(_367_),
    .B1(_357_),
    .X(_283_));
 sky130_fd_sc_hd__a21o_1 _728_ (.A1(_343_),
    .A2(_374_),
    .B1(net41),
    .X(_284_));
 sky130_fd_sc_hd__o211ai_1 _729_ (.A1(net26),
    .A2(_283_),
    .B1(_284_),
    .C1(_347_),
    .Y(_285_));
 sky130_fd_sc_hd__o221a_1 _730_ (.A1(_373_),
    .A2(_019_),
    .B1(_075_),
    .B2(_353_),
    .C1(net26),
    .X(_286_));
 sky130_fd_sc_hd__a211o_1 _731_ (.A1(net55),
    .A2(net19),
    .B1(_349_),
    .C1(_371_),
    .X(_287_));
 sky130_fd_sc_hd__o211a_1 _732_ (.A1(net45),
    .A2(_197_),
    .B1(_287_),
    .C1(net35),
    .X(_288_));
 sky130_fd_sc_hd__o31a_1 _733_ (.A1(_032_),
    .A2(_286_),
    .A3(_288_),
    .B1(_285_),
    .X(_289_));
 sky130_fd_sc_hd__nand2_1 _734_ (.A(_372_),
    .B(_028_),
    .Y(_290_));
 sky130_fd_sc_hd__a21oi_1 _735_ (.A1(_001_),
    .A2(_023_),
    .B1(_129_),
    .Y(_291_));
 sky130_fd_sc_hd__a211o_1 _736_ (.A1(net38),
    .A2(_290_),
    .B1(_291_),
    .C1(_052_),
    .X(_292_));
 sky130_fd_sc_hd__nand2_1 _737_ (.A(_372_),
    .B(_076_),
    .Y(_293_));
 sky130_fd_sc_hd__or2_1 _738_ (.A(net27),
    .B(_384_),
    .X(_294_));
 sky130_fd_sc_hd__a31o_1 _739_ (.A1(net20),
    .A2(_111_),
    .A3(_293_),
    .B1(_294_),
    .X(_295_));
 sky130_fd_sc_hd__or4_1 _740_ (.A(net36),
    .B(_351_),
    .C(_384_),
    .D(_260_),
    .X(_296_));
 sky130_fd_sc_hd__a21o_1 _741_ (.A1(_295_),
    .A2(_296_),
    .B1(net21),
    .X(_297_));
 sky130_fd_sc_hd__and3_1 _742_ (.A(_289_),
    .B(_292_),
    .C(_297_),
    .X(_298_));
 sky130_fd_sc_hd__or3_1 _743_ (.A(net35),
    .B(_069_),
    .C(_092_),
    .X(_299_));
 sky130_fd_sc_hd__or3_1 _744_ (.A(net35),
    .B(net25),
    .C(_026_),
    .X(_300_));
 sky130_fd_sc_hd__a31o_1 _745_ (.A1(_295_),
    .A2(_299_),
    .A3(_300_),
    .B1(net21),
    .X(_301_));
 sky130_fd_sc_hd__and3_1 _746_ (.A(net30),
    .B(_289_),
    .C(_292_),
    .X(_302_));
 sky130_fd_sc_hd__o2bb2a_1 _747_ (.A1_N(_301_),
    .A2_N(_302_),
    .B1(net30),
    .B2(_298_),
    .X(net3));
 sky130_fd_sc_hd__or3b_1 _748_ (.A(_161_),
    .B(_294_),
    .C_N(_179_),
    .X(_303_));
 sky130_fd_sc_hd__a31o_1 _749_ (.A1(_016_),
    .A2(_023_),
    .A3(_063_),
    .B1(net42),
    .X(_304_));
 sky130_fd_sc_hd__o2111a_1 _750_ (.A1(_374_),
    .A2(_090_),
    .B1(_035_),
    .C1(_337_),
    .D1(net43),
    .X(_305_));
 sky130_fd_sc_hd__a311o_1 _751_ (.A1(net33),
    .A2(_303_),
    .A3(_304_),
    .B1(_305_),
    .C1(_331_),
    .X(_306_));
 sky130_fd_sc_hd__a211o_1 _752_ (.A1(_360_),
    .A2(_372_),
    .B1(_082_),
    .C1(net42),
    .X(_307_));
 sky130_fd_sc_hd__nand2_1 _753_ (.A(net42),
    .B(_065_),
    .Y(_308_));
 sky130_fd_sc_hd__a31oi_1 _754_ (.A1(net33),
    .A2(_307_),
    .A3(_308_),
    .B1(\tcount[6] ),
    .Y(_309_));
 sky130_fd_sc_hd__a21o_1 _755_ (.A1(_368_),
    .A2(net20),
    .B1(net53),
    .X(_310_));
 sky130_fd_sc_hd__o311a_1 _756_ (.A1(net24),
    .A2(_367_),
    .A3(_036_),
    .B1(_086_),
    .C1(net39),
    .X(_311_));
 sky130_fd_sc_hd__a311o_1 _757_ (.A1(net29),
    .A2(_377_),
    .A3(_310_),
    .B1(_311_),
    .C1(net33),
    .X(_312_));
 sky130_fd_sc_hd__nand2_1 _758_ (.A(_309_),
    .B(_312_),
    .Y(_313_));
 sky130_fd_sc_hd__o21ai_1 _759_ (.A1(_184_),
    .A2(_311_),
    .B1(_309_),
    .Y(_314_));
 sky130_fd_sc_hd__a21oi_1 _760_ (.A1(_306_),
    .A2(_314_),
    .B1(net31),
    .Y(_315_));
 sky130_fd_sc_hd__a31o_1 _761_ (.A1(net31),
    .A2(_306_),
    .A3(_313_),
    .B1(_315_),
    .X(net4));
 sky130_fd_sc_hd__a211o_1 _762_ (.A1(net68),
    .A2(_384_),
    .B1(_134_),
    .C1(net40),
    .X(_316_));
 sky130_fd_sc_hd__o31ai_1 _763_ (.A1(_349_),
    .A2(_363_),
    .A3(_134_),
    .B1(net40),
    .Y(_317_));
 sky130_fd_sc_hd__a31o_1 _764_ (.A1(_337_),
    .A2(net40),
    .A3(_091_),
    .B1(_331_),
    .X(_318_));
 sky130_fd_sc_hd__a31o_1 _765_ (.A1(net34),
    .A2(_316_),
    .A3(_317_),
    .B1(_318_),
    .X(_319_));
 sky130_fd_sc_hd__a22o_1 _766_ (.A1(net49),
    .A2(_359_),
    .B1(_076_),
    .B2(net58),
    .X(_320_));
 sky130_fd_sc_hd__and2_1 _767_ (.A(net27),
    .B(_320_),
    .X(_321_));
 sky130_fd_sc_hd__a21oi_1 _768_ (.A1(net40),
    .A2(_350_),
    .B1(_134_),
    .Y(_322_));
 sky130_fd_sc_hd__a31o_1 _769_ (.A1(net40),
    .A2(net49),
    .A3(_359_),
    .B1(_389_),
    .X(_323_));
 sky130_fd_sc_hd__o221a_1 _770_ (.A1(_052_),
    .A2(_321_),
    .B1(_322_),
    .B2(_323_),
    .C1(_319_),
    .X(_324_));
 sky130_fd_sc_hd__or2_1 _771_ (.A(net43),
    .B(_179_),
    .X(_325_));
 sky130_fd_sc_hd__and2_1 _772_ (.A(net31),
    .B(_325_),
    .X(_326_));
 sky130_fd_sc_hd__mux2_1 _773_ (.A0(_341_),
    .A1(_326_),
    .S(_324_),
    .X(net5));
 sky130_fd_sc_hd__a22o_1 _774_ (.A1(_051_),
    .A2(_183_),
    .B1(_284_),
    .B2(_145_),
    .X(_327_));
 sky130_fd_sc_hd__or2_1 _775_ (.A(_347_),
    .B(_327_),
    .X(_328_));
 sky130_fd_sc_hd__o21a_1 _776_ (.A1(net33),
    .A2(_325_),
    .B1(net31),
    .X(_329_));
 sky130_fd_sc_hd__mux2_1 _777_ (.A0(_329_),
    .A1(_341_),
    .S(_328_),
    .X(net6));
 sky130_fd_sc_hd__a32oi_2 _778_ (.A1(_388_),
    .A2(_145_),
    .A3(_325_),
    .B1(_284_),
    .B2(_031_),
    .Y(_330_));
 sky130_fd_sc_hd__or3_1 _779_ (.A(\tcount[6] ),
    .B(net33),
    .C(_325_),
    .X(_332_));
 sky130_fd_sc_hd__a21oi_1 _780_ (.A1(_330_),
    .A2(_332_),
    .B1(net31),
    .Y(_333_));
 sky130_fd_sc_hd__a21oi_1 _781_ (.A1(net31),
    .A2(_330_),
    .B1(_333_),
    .Y(net7));
 sky130_fd_sc_hd__and2_1 _782_ (.A(net32),
    .B(_332_),
    .X(net8));
 sky130_fd_sc_hd__nor2_1 _783_ (.A(_090_),
    .B(_128_),
    .Y(_003_));
 sky130_fd_sc_hd__nand2_1 _784_ (.A(net43),
    .B(_128_),
    .Y(_334_));
 sky130_fd_sc_hd__and2_1 _785_ (.A(_129_),
    .B(_334_),
    .X(_004_));
 sky130_fd_sc_hd__xnor2_1 _786_ (.A(net34),
    .B(_334_),
    .Y(_005_));
 sky130_fd_sc_hd__or2_1 _787_ (.A(_032_),
    .B(_334_),
    .X(_335_));
 sky130_fd_sc_hd__a31o_1 _788_ (.A1(net34),
    .A2(net43),
    .A3(_128_),
    .B1(\tcount[6] ),
    .X(_336_));
 sky130_fd_sc_hd__and2_1 _789_ (.A(_335_),
    .B(_336_),
    .X(_006_));
 sky130_fd_sc_hd__xnor2_1 _790_ (.A(net32),
    .B(_335_),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _791_ (.A(net1),
    .Y(_009_));
 sky130_fd_sc_hd__inv_2 _792_ (.A(net1),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _793_ (.A(net1),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _794_ (.A(net1),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _795_ (.A(net1),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _796_ (.A(net1),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _797_ (.A(net1),
    .Y(_015_));
 sky130_fd_sc_hd__dfrtp_1 _798_ (.CLK(clknet_1_0__leaf_clk),
    .D(_000_),
    .RESET_B(_008_),
    .Q(\tcount[0] ));
 sky130_fd_sc_hd__dfrtp_1 _799_ (.CLK(clknet_1_0__leaf_clk),
    .D(net19),
    .RESET_B(_009_),
    .Q(\tcount[1] ));
 sky130_fd_sc_hd__dfrtp_2 _800_ (.CLK(clknet_1_0__leaf_clk),
    .D(_002_),
    .RESET_B(_010_),
    .Q(\tcount[2] ));
 sky130_fd_sc_hd__dfrtp_1 _801_ (.CLK(clknet_1_0__leaf_clk),
    .D(_003_),
    .RESET_B(_011_),
    .Q(\tcount[3] ));
 sky130_fd_sc_hd__dfrtp_1 _802_ (.CLK(clknet_1_1__leaf_clk),
    .D(_004_),
    .RESET_B(_012_),
    .Q(\tcount[4] ));
 sky130_fd_sc_hd__dfrtp_1 _803_ (.CLK(clknet_1_1__leaf_clk),
    .D(_005_),
    .RESET_B(_013_),
    .Q(\tcount[5] ));
 sky130_fd_sc_hd__dfrtp_4 _804_ (.CLK(clknet_1_1__leaf_clk),
    .D(_006_),
    .RESET_B(_014_),
    .Q(\tcount[6] ));
 sky130_fd_sc_hd__dfrtp_1 _805_ (.CLK(clknet_1_1__leaf_clk),
    .D(_007_),
    .RESET_B(_015_),
    .Q(\tcount[7] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_160 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(rst),
    .X(net1));
 sky130_fd_sc_hd__buf_2 output2 (.A(net2),
    .X(sine_out[0]));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(sine_out[10]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(sine_out[11]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(sine_out[12]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(sine_out[13]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(sine_out[14]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(sine_out[15]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(sine_out[1]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(sine_out[2]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(sine_out[3]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(sine_out[4]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(sine_out[5]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(sine_out[6]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(sine_out[7]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(sine_out[8]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(sine_out[9]));
 sky130_fd_sc_hd__buf_1 max_cap18 (.A(_047_),
    .X(net18));
 sky130_fd_sc_hd__buf_2 fanout19 (.A(_001_),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 fanout20 (.A(_037_),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 fanout21 (.A(_389_),
    .X(net21));
 sky130_fd_sc_hd__buf_2 fanout22 (.A(_360_),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 fanout23 (.A(_346_),
    .X(net23));
 sky130_fd_sc_hd__buf_2 fanout24 (.A(net25),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 fanout25 (.A(_339_),
    .X(net25));
 sky130_fd_sc_hd__buf_2 fanout26 (.A(net29),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__buf_2 fanout29 (.A(_338_),
    .X(net29));
 sky130_fd_sc_hd__buf_2 fanout30 (.A(net32),
    .X(net30));
 sky130_fd_sc_hd__buf_2 fanout31 (.A(net32),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 fanout32 (.A(\tcount[7] ),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 fanout33 (.A(net34),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 fanout34 (.A(\tcount[5] ),
    .X(net34));
 sky130_fd_sc_hd__buf_2 fanout35 (.A(net39),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 fanout36 (.A(net39),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout39 (.A(net44),
    .X(net39));
 sky130_fd_sc_hd__buf_2 fanout40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(net44),
    .X(net41));
 sky130_fd_sc_hd__buf_2 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout44 (.A(\tcount[4] ),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(net49),
    .X(net46));
 sky130_fd_sc_hd__buf_2 fanout47 (.A(net49),
    .X(net47));
 sky130_fd_sc_hd__buf_2 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__buf_2 fanout49 (.A(net54),
    .X(net49));
 sky130_fd_sc_hd__buf_2 fanout50 (.A(net54),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net54),
    .X(net51));
 sky130_fd_sc_hd__buf_2 fanout52 (.A(net54),
    .X(net52));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 fanout54 (.A(\tcount[3] ),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__buf_2 fanout56 (.A(\tcount[2] ),
    .X(net56));
 sky130_fd_sc_hd__buf_4 fanout57 (.A(\tcount[2] ),
    .X(net57));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout58 (.A(\tcount[2] ),
    .X(net58));
 sky130_fd_sc_hd__buf_2 fanout59 (.A(net61),
    .X(net59));
 sky130_fd_sc_hd__buf_2 fanout60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 fanout61 (.A(\tcount[2] ),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(net64),
    .X(net62));
 sky130_fd_sc_hd__buf_4 fanout63 (.A(net64),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 fanout64 (.A(\tcount[1] ),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 fanout65 (.A(net66),
    .X(net65));
 sky130_fd_sc_hd__buf_2 fanout66 (.A(\tcount[1] ),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 fanout67 (.A(net70),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 fanout68 (.A(net70),
    .X(net68));
 sky130_fd_sc_hd__buf_1 fanout69 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__buf_2 fanout70 (.A(\tcount[0] ),
    .X(net70));
 sky130_fd_sc_hd__buf_4 fanout71 (.A(net72),
    .X(net71));
 sky130_fd_sc_hd__buf_2 fanout72 (.A(\tcount[0] ),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_181 ();
endmodule
