module counter_8bit (clk,
    rst,
    sine_out);
 input clk;
 input rst;
 output [15:0] sine_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire \tcount[0] ;
 wire \tcount[1] ;
 wire \tcount[2] ;
 wire \tcount[3] ;
 wire \tcount[4] ;
 wire \tcount[5] ;
 wire \tcount[6] ;
 wire \tcount[7] ;

 sky130_fd_sc_hd__inv_2 _391_ (.A(\tcount[0] ),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _392_ (.A(\tcount[6] ),
    .Y(_331_));
 sky130_fd_sc_hd__inv_2 _393_ (.A(\tcount[5] ),
    .Y(_337_));
 sky130_fd_sc_hd__inv_2 _394_ (.A(\tcount[4] ),
    .Y(_338_));
 sky130_fd_sc_hd__inv_2 _395_ (.A(\tcount[3] ),
    .Y(_339_));
 sky130_fd_sc_hd__inv_2 _396_ (.A(\tcount[1] ),
    .Y(_340_));
 sky130_fd_sc_hd__inv_2 _397_ (.A(\tcount[7] ),
    .Y(_341_));
 sky130_fd_sc_hd__inv_2 _398_ (.A(rst),
    .Y(_008_));
 sky130_fd_sc_hd__nor2_2 _399_ (.A(\tcount[0] ),
    .B(\tcount[1] ),
    .Y(_342_));
 sky130_fd_sc_hd__or2_2 _400_ (.A(\tcount[0] ),
    .B(\tcount[1] ),
    .X(_343_));
 sky130_fd_sc_hd__and2_2 _401_ (.A(\tcount[0] ),
    .B(\tcount[1] ),
    .X(_344_));
 sky130_fd_sc_hd__nand2_2 _402_ (.A(\tcount[0] ),
    .B(\tcount[1] ),
    .Y(_345_));
 sky130_fd_sc_hd__xnor2_2 _403_ (.A(\tcount[0] ),
    .B(\tcount[1] ),
    .Y(_346_));
 sky130_fd_sc_hd__inv_2 _404_ (.A(_346_),
    .Y(_001_));
 sky130_fd_sc_hd__nor2_2 _405_ (.A(_331_),
    .B(\tcount[5] ),
    .Y(_347_));
 sky130_fd_sc_hd__nand2_2 _406_ (.A(\tcount[6] ),
    .B(_337_),
    .Y(_348_));
 sky130_fd_sc_hd__nor2_2 _407_ (.A(\tcount[2] ),
    .B(\tcount[1] ),
    .Y(_349_));
 sky130_fd_sc_hd__or2_2 _408_ (.A(\tcount[2] ),
    .B(\tcount[1] ),
    .X(_350_));
 sky130_fd_sc_hd__and2b_2 _409_ (.A_N(\tcount[0] ),
    .B(\tcount[2] ),
    .X(_351_));
 sky130_fd_sc_hd__nand2b_2 _410_ (.A_N(\tcount[0] ),
    .B(\tcount[2] ),
    .Y(_352_));
 sky130_fd_sc_hd__and2b_2 _411_ (.A_N(\tcount[2] ),
    .B(\tcount[1] ),
    .X(_353_));
 sky130_fd_sc_hd__nand2b_2 _412_ (.A_N(\tcount[2] ),
    .B(\tcount[1] ),
    .Y(_354_));
 sky130_fd_sc_hd__and2_2 _413_ (.A(\tcount[0] ),
    .B(\tcount[2] ),
    .X(_355_));
 sky130_fd_sc_hd__nand2_2 _414_ (.A(\tcount[0] ),
    .B(\tcount[2] ),
    .Y(_356_));
 sky130_fd_sc_hd__nand2b_2 _415_ (.A_N(\tcount[1] ),
    .B(\tcount[3] ),
    .Y(_357_));
 sky130_fd_sc_hd__nand2b_2 _416_ (.A_N(\tcount[2] ),
    .B(\tcount[3] ),
    .Y(_358_));
 sky130_fd_sc_hd__nand2_2 _417_ (.A(\tcount[2] ),
    .B(\tcount[1] ),
    .Y(_359_));
 sky130_fd_sc_hd__xnor2_2 _418_ (.A(\tcount[2] ),
    .B(\tcount[1] ),
    .Y(_360_));
 sky130_fd_sc_hd__o21ai_2 _419_ (.A1(\tcount[0] ),
    .A2(\tcount[1] ),
    .B1(\tcount[3] ),
    .Y(_361_));
 sky130_fd_sc_hd__inv_2 _420_ (.A(_361_),
    .Y(_362_));
 sky130_fd_sc_hd__nor2_2 _421_ (.A(\tcount[0] ),
    .B(\tcount[2] ),
    .Y(_363_));
 sky130_fd_sc_hd__o21ai_2 _422_ (.A1(\tcount[0] ),
    .A2(\tcount[2] ),
    .B1(\tcount[3] ),
    .Y(_364_));
 sky130_fd_sc_hd__nor3_2 _423_ (.A(_000_),
    .B(_339_),
    .C(_360_),
    .Y(_365_));
 sky130_fd_sc_hd__nor2_2 _424_ (.A(\tcount[2] ),
    .B(_346_),
    .Y(_366_));
 sky130_fd_sc_hd__and2b_2 _425_ (.A_N(\tcount[1] ),
    .B(\tcount[2] ),
    .X(_367_));
 sky130_fd_sc_hd__or3b_2 _426_ (.A(\tcount[0] ),
    .B(\tcount[1] ),
    .C_N(\tcount[2] ),
    .X(_368_));
 sky130_fd_sc_hd__o211ai_2 _427_ (.A1(\tcount[2] ),
    .A2(_346_),
    .B1(_368_),
    .C1(_339_),
    .Y(_369_));
 sky130_fd_sc_hd__nand2_2 _428_ (.A(\tcount[4] ),
    .B(_369_),
    .Y(_370_));
 sky130_fd_sc_hd__and2b_2 _429_ (.A_N(\tcount[2] ),
    .B(\tcount[0] ),
    .X(_371_));
 sky130_fd_sc_hd__nand2b_2 _430_ (.A_N(\tcount[2] ),
    .B(\tcount[0] ),
    .Y(_372_));
 sky130_fd_sc_hd__and2_2 _431_ (.A(\tcount[2] ),
    .B(_346_),
    .X(_373_));
 sky130_fd_sc_hd__and2_2 _432_ (.A(\tcount[3] ),
    .B(\tcount[2] ),
    .X(_374_));
 sky130_fd_sc_hd__nand2_2 _433_ (.A(\tcount[3] ),
    .B(\tcount[2] ),
    .Y(_375_));
 sky130_fd_sc_hd__nand2_2 _434_ (.A(\tcount[3] ),
    .B(_354_),
    .Y(_376_));
 sky130_fd_sc_hd__a211o_2 _435_ (.A1(\tcount[2] ),
    .A2(_346_),
    .B1(_353_),
    .C1(_339_),
    .X(_377_));
 sky130_fd_sc_hd__nor2_2 _436_ (.A(_371_),
    .B(_377_),
    .Y(_378_));
 sky130_fd_sc_hd__nor3_2 _437_ (.A(\tcount[0] ),
    .B(\tcount[3] ),
    .C(\tcount[1] ),
    .Y(_379_));
 sky130_fd_sc_hd__nor3b_2 _438_ (.A(\tcount[3] ),
    .B(\tcount[1] ),
    .C_N(\tcount[2] ),
    .Y(_380_));
 sky130_fd_sc_hd__nand2_2 _439_ (.A(_339_),
    .B(_367_),
    .Y(_381_));
 sky130_fd_sc_hd__or4_2 _440_ (.A(\tcount[4] ),
    .B(_378_),
    .C(_379_),
    .D(_380_),
    .X(_382_));
 sky130_fd_sc_hd__o21ai_2 _441_ (.A1(_365_),
    .A2(_370_),
    .B1(_382_),
    .Y(_383_));
 sky130_fd_sc_hd__and3b_2 _442_ (.A_N(\tcount[3] ),
    .B(\tcount[2] ),
    .C(\tcount[1] ),
    .X(_384_));
 sky130_fd_sc_hd__nor2_2 _443_ (.A(\tcount[4] ),
    .B(_384_),
    .Y(_385_));
 sky130_fd_sc_hd__nor2_2 _444_ (.A(\tcount[0] ),
    .B(\tcount[4] ),
    .Y(_386_));
 sky130_fd_sc_hd__o22a_2 _445_ (.A1(_360_),
    .A2(_361_),
    .B1(_385_),
    .B2(_386_),
    .X(_387_));
 sky130_fd_sc_hd__nor2_2 _446_ (.A(\tcount[6] ),
    .B(\tcount[5] ),
    .Y(_388_));
 sky130_fd_sc_hd__or2_2 _447_ (.A(\tcount[6] ),
    .B(\tcount[5] ),
    .X(_389_));
 sky130_fd_sc_hd__a21bo_2 _448_ (.A1(\tcount[0] ),
    .A2(\tcount[1] ),
    .B1_N(\tcount[2] ),
    .X(_390_));
 sky130_fd_sc_hd__nand2_2 _449_ (.A(_339_),
    .B(_390_),
    .Y(_016_));
 sky130_fd_sc_hd__a31o_2 _450_ (.A1(\tcount[4] ),
    .A2(_375_),
    .A3(_016_),
    .B1(_389_),
    .X(_017_));
 sky130_fd_sc_hd__o21ba_2 _451_ (.A1(\tcount[2] ),
    .A2(\tcount[1] ),
    .B1_N(\tcount[3] ),
    .X(_018_));
 sky130_fd_sc_hd__o21bai_2 _452_ (.A1(\tcount[2] ),
    .A2(\tcount[1] ),
    .B1_N(\tcount[3] ),
    .Y(_019_));
 sky130_fd_sc_hd__nor2_2 _453_ (.A(_001_),
    .B(_019_),
    .Y(_020_));
 sky130_fd_sc_hd__and2b_2 _454_ (.A_N(\tcount[1] ),
    .B(\tcount[0] ),
    .X(_021_));
 sky130_fd_sc_hd__nand2b_2 _455_ (.A_N(\tcount[1] ),
    .B(\tcount[0] ),
    .Y(_022_));
 sky130_fd_sc_hd__nand2_2 _456_ (.A(\tcount[3] ),
    .B(_355_),
    .Y(_023_));
 sky130_fd_sc_hd__nor2_2 _457_ (.A(_375_),
    .B(_022_),
    .Y(_024_));
 sky130_fd_sc_hd__nor2_2 _458_ (.A(_351_),
    .B(_371_),
    .Y(_025_));
 sky130_fd_sc_hd__xor2_2 _459_ (.A(\tcount[0] ),
    .B(\tcount[2] ),
    .X(_026_));
 sky130_fd_sc_hd__or2_2 _460_ (.A(\tcount[1] ),
    .B(_026_),
    .X(_027_));
 sky130_fd_sc_hd__nor2_2 _461_ (.A(\tcount[3] ),
    .B(_353_),
    .Y(_028_));
 sky130_fd_sc_hd__a21oi_2 _462_ (.A1(_339_),
    .A2(_354_),
    .B1(\tcount[4] ),
    .Y(_029_));
 sky130_fd_sc_hd__nand2_2 _463_ (.A(_027_),
    .B(_029_),
    .Y(_030_));
 sky130_fd_sc_hd__nor2_2 _464_ (.A(_331_),
    .B(_337_),
    .Y(_031_));
 sky130_fd_sc_hd__nand2_2 _465_ (.A(\tcount[6] ),
    .B(\tcount[5] ),
    .Y(_032_));
 sky130_fd_sc_hd__o41a_2 _466_ (.A1(_338_),
    .A2(_366_),
    .A3(_020_),
    .A4(_024_),
    .B1(_031_),
    .X(_033_));
 sky130_fd_sc_hd__a2bb2o_2 _467_ (.A1_N(_387_),
    .A2_N(_017_),
    .B1(_030_),
    .B2(_033_),
    .X(_034_));
 sky130_fd_sc_hd__or3_2 _468_ (.A(\tcount[0] ),
    .B(\tcount[2] ),
    .C(\tcount[1] ),
    .X(_035_));
 sky130_fd_sc_hd__and3b_2 _469_ (.A_N(\tcount[2] ),
    .B(\tcount[1] ),
    .C(\tcount[0] ),
    .X(_036_));
 sky130_fd_sc_hd__nand3b_2 _470_ (.A_N(\tcount[2] ),
    .B(\tcount[1] ),
    .C(\tcount[0] ),
    .Y(_037_));
 sky130_fd_sc_hd__nand2_2 _471_ (.A(_390_),
    .B(_037_),
    .Y(_002_));
 sky130_fd_sc_hd__and3_2 _472_ (.A(_390_),
    .B(_035_),
    .C(_037_),
    .X(_038_));
 sky130_fd_sc_hd__nand2_2 _473_ (.A(\tcount[3] ),
    .B(\tcount[1] ),
    .Y(_039_));
 sky130_fd_sc_hd__nand2_2 _474_ (.A(_375_),
    .B(_039_),
    .Y(_040_));
 sky130_fd_sc_hd__a21bo_2 _475_ (.A1(\tcount[0] ),
    .A2(\tcount[1] ),
    .B1_N(\tcount[3] ),
    .X(_041_));
 sky130_fd_sc_hd__nand2_2 _476_ (.A(\tcount[3] ),
    .B(_372_),
    .Y(_042_));
 sky130_fd_sc_hd__a21oi_2 _477_ (.A1(_001_),
    .A2(_040_),
    .B1(_038_),
    .Y(_043_));
 sky130_fd_sc_hd__and3_2 _478_ (.A(\tcount[3] ),
    .B(\tcount[1] ),
    .C(_363_),
    .X(_044_));
 sky130_fd_sc_hd__nor3b_2 _479_ (.A(\tcount[2] ),
    .B(\tcount[1] ),
    .C_N(\tcount[0] ),
    .Y(_045_));
 sky130_fd_sc_hd__nor2_2 _480_ (.A(\tcount[3] ),
    .B(_045_),
    .Y(_046_));
 sky130_fd_sc_hd__nor3_2 _481_ (.A(\tcount[3] ),
    .B(_351_),
    .C(_045_),
    .Y(_047_));
 sky130_fd_sc_hd__and2_2 _482_ (.A(_359_),
    .B(_047_),
    .X(_048_));
 sky130_fd_sc_hd__a21o_2 _483_ (.A1(\tcount[2] ),
    .A2(_346_),
    .B1(_339_),
    .X(_049_));
 sky130_fd_sc_hd__or3b_2 _484_ (.A(_338_),
    .B(_048_),
    .C_N(_049_),
    .X(_050_));
 sky130_fd_sc_hd__nor2_2 _485_ (.A(\tcount[6] ),
    .B(_337_),
    .Y(_051_));
 sky130_fd_sc_hd__nand2_2 _486_ (.A(_331_),
    .B(\tcount[5] ),
    .Y(_052_));
 sky130_fd_sc_hd__o311a_2 _487_ (.A1(\tcount[4] ),
    .A2(_043_),
    .A3(_044_),
    .B1(_050_),
    .C1(_051_),
    .X(_053_));
 sky130_fd_sc_hd__a211o_2 _488_ (.A1(_347_),
    .A2(_383_),
    .B1(_034_),
    .C1(_053_),
    .X(sine_out[0]));
 sky130_fd_sc_hd__a221oi_2 _489_ (.A1(_000_),
    .A2(_380_),
    .B1(_038_),
    .B2(\tcount[3] ),
    .C1(_032_),
    .Y(_054_));
 sky130_fd_sc_hd__a32o_2 _490_ (.A1(_345_),
    .A2(_018_),
    .A3(_025_),
    .B1(_036_),
    .B2(\tcount[3] ),
    .X(_055_));
 sky130_fd_sc_hd__nor2_2 _491_ (.A(_342_),
    .B(_390_),
    .Y(_056_));
 sky130_fd_sc_hd__nand2_2 _492_ (.A(\tcount[2] ),
    .B(_001_),
    .Y(_057_));
 sky130_fd_sc_hd__nor2_2 _493_ (.A(_349_),
    .B(_042_),
    .Y(_058_));
 sky130_fd_sc_hd__and2_2 _494_ (.A(_339_),
    .B(_360_),
    .X(_059_));
 sky130_fd_sc_hd__and3_2 _495_ (.A(_339_),
    .B(_360_),
    .C(_022_),
    .X(_060_));
 sky130_fd_sc_hd__a31oi_2 _496_ (.A1(_372_),
    .A2(_040_),
    .A3(_057_),
    .B1(_060_),
    .Y(_061_));
 sky130_fd_sc_hd__a221o_2 _497_ (.A1(_347_),
    .A2(_055_),
    .B1(_061_),
    .B2(_051_),
    .C1(_054_),
    .X(_062_));
 sky130_fd_sc_hd__nand2_2 _498_ (.A(\tcount[3] ),
    .B(_360_),
    .Y(_063_));
 sky130_fd_sc_hd__nor2_2 _499_ (.A(\tcount[3] ),
    .B(\tcount[2] ),
    .Y(_064_));
 sky130_fd_sc_hd__or2_2 _500_ (.A(\tcount[3] ),
    .B(\tcount[2] ),
    .X(_065_));
 sky130_fd_sc_hd__nand2b_2 _501_ (.A_N(\tcount[3] ),
    .B(\tcount[0] ),
    .Y(_066_));
 sky130_fd_sc_hd__nor2_2 _502_ (.A(_345_),
    .B(_065_),
    .Y(_067_));
 sky130_fd_sc_hd__a31o_2 _503_ (.A1(\tcount[0] ),
    .A2(\tcount[3] ),
    .A3(_360_),
    .B1(_067_),
    .X(_068_));
 sky130_fd_sc_hd__o21ba_2 _504_ (.A1(\tcount[2] ),
    .A2(\tcount[1] ),
    .B1_N(\tcount[0] ),
    .X(_069_));
 sky130_fd_sc_hd__o21bai_2 _505_ (.A1(\tcount[2] ),
    .A2(\tcount[1] ),
    .B1_N(\tcount[0] ),
    .Y(_070_));
 sky130_fd_sc_hd__nand2_2 _506_ (.A(\tcount[3] ),
    .B(_070_),
    .Y(_071_));
 sky130_fd_sc_hd__nand2_2 _507_ (.A(\tcount[1] ),
    .B(_026_),
    .Y(_072_));
 sky130_fd_sc_hd__a21bo_2 _508_ (.A1(_339_),
    .A2(_072_),
    .B1_N(_071_),
    .X(_073_));
 sky130_fd_sc_hd__a21oi_2 _509_ (.A1(\tcount[2] ),
    .A2(_001_),
    .B1(_364_),
    .Y(_074_));
 sky130_fd_sc_hd__a21o_2 _510_ (.A1(\tcount[2] ),
    .A2(_001_),
    .B1(_364_),
    .X(_075_));
 sky130_fd_sc_hd__o21ba_2 _511_ (.A1(\tcount[0] ),
    .A2(\tcount[1] ),
    .B1_N(\tcount[3] ),
    .X(_076_));
 sky130_fd_sc_hd__nand2_2 _512_ (.A(_360_),
    .B(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__a21oi_2 _513_ (.A1(_075_),
    .A2(_077_),
    .B1(_348_),
    .Y(_078_));
 sky130_fd_sc_hd__a221o_2 _514_ (.A1(_051_),
    .A2(_068_),
    .B1(_073_),
    .B2(_031_),
    .C1(_338_),
    .X(_079_));
 sky130_fd_sc_hd__o22a_2 _515_ (.A1(\tcount[4] ),
    .A2(_062_),
    .B1(_078_),
    .B2(_079_),
    .X(_080_));
 sky130_fd_sc_hd__a21o_2 _516_ (.A1(\tcount[1] ),
    .A2(_351_),
    .B1(_364_),
    .X(_081_));
 sky130_fd_sc_hd__and3b_2 _517_ (.A_N(\tcount[3] ),
    .B(\tcount[2] ),
    .C(\tcount[0] ),
    .X(_082_));
 sky130_fd_sc_hd__nor2_2 _518_ (.A(\tcount[4] ),
    .B(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__o211a_2 _519_ (.A1(\tcount[3] ),
    .A2(_021_),
    .B1(_376_),
    .C1(\tcount[4] ),
    .X(_084_));
 sky130_fd_sc_hd__a211oi_2 _520_ (.A1(_081_),
    .A2(_083_),
    .B1(_084_),
    .C1(_389_),
    .Y(_085_));
 sky130_fd_sc_hd__or3_2 _521_ (.A(\tcount[3] ),
    .B(_360_),
    .C(_021_),
    .X(_086_));
 sky130_fd_sc_hd__nor2_2 _522_ (.A(_349_),
    .B(_364_),
    .Y(_087_));
 sky130_fd_sc_hd__o311a_2 _523_ (.A1(_349_),
    .A2(_355_),
    .A3(_364_),
    .B1(_086_),
    .C1(_338_),
    .X(_088_));
 sky130_fd_sc_hd__and3_2 _524_ (.A(\tcount[0] ),
    .B(\tcount[2] ),
    .C(\tcount[1] ),
    .X(_089_));
 sky130_fd_sc_hd__nor2_2 _525_ (.A(\tcount[3] ),
    .B(_089_),
    .Y(_090_));
 sky130_fd_sc_hd__a31o_2 _526_ (.A1(\tcount[0] ),
    .A2(\tcount[2] ),
    .A3(\tcount[1] ),
    .B1(\tcount[3] ),
    .X(_091_));
 sky130_fd_sc_hd__or2_2 _527_ (.A(_045_),
    .B(_091_),
    .X(_092_));
 sky130_fd_sc_hd__o31a_2 _528_ (.A1(_339_),
    .A2(_351_),
    .A3(_021_),
    .B1(\tcount[4] ),
    .X(_093_));
 sky130_fd_sc_hd__o21a_2 _529_ (.A1(_069_),
    .A2(_092_),
    .B1(_093_),
    .X(_094_));
 sky130_fd_sc_hd__a311o_2 _530_ (.A1(\tcount[3] ),
    .A2(_340_),
    .A3(_363_),
    .B1(_380_),
    .C1(_344_),
    .X(_095_));
 sky130_fd_sc_hd__nor2_2 _531_ (.A(_357_),
    .B(_371_),
    .Y(_096_));
 sky130_fd_sc_hd__o211a_2 _532_ (.A1(_344_),
    .A2(_026_),
    .B1(_039_),
    .C1(\tcount[4] ),
    .X(_097_));
 sky130_fd_sc_hd__a211o_2 _533_ (.A1(_338_),
    .A2(_095_),
    .B1(_097_),
    .C1(_052_),
    .X(_098_));
 sky130_fd_sc_hd__o311a_2 _534_ (.A1(_032_),
    .A2(_088_),
    .A3(_094_),
    .B1(_098_),
    .C1(\tcount[7] ),
    .X(_099_));
 sky130_fd_sc_hd__inv_2 _535_ (.A(_099_),
    .Y(_100_));
 sky130_fd_sc_hd__and3_2 _536_ (.A(\tcount[3] ),
    .B(_027_),
    .C(_072_),
    .X(_101_));
 sky130_fd_sc_hd__a211o_2 _537_ (.A1(\tcount[0] ),
    .A2(_380_),
    .B1(_101_),
    .C1(\tcount[4] ),
    .X(_102_));
 sky130_fd_sc_hd__a21o_2 _538_ (.A1(\tcount[3] ),
    .A2(_349_),
    .B1(_338_),
    .X(_103_));
 sky130_fd_sc_hd__a21o_2 _539_ (.A1(_026_),
    .A2(_028_),
    .B1(_103_),
    .X(_104_));
 sky130_fd_sc_hd__nand2_2 _540_ (.A(_385_),
    .B(_066_),
    .Y(_105_));
 sky130_fd_sc_hd__a21o_2 _541_ (.A1(_000_),
    .A2(\tcount[1] ),
    .B1(_338_),
    .X(_106_));
 sky130_fd_sc_hd__nand2_2 _542_ (.A(_375_),
    .B(_065_),
    .Y(_107_));
 sky130_fd_sc_hd__a31o_2 _543_ (.A1(_375_),
    .A2(_022_),
    .A3(_065_),
    .B1(_106_),
    .X(_108_));
 sky130_fd_sc_hd__o211a_2 _544_ (.A1(_101_),
    .A2(_105_),
    .B1(_108_),
    .C1(_347_),
    .X(_109_));
 sky130_fd_sc_hd__a31o_2 _545_ (.A1(_388_),
    .A2(_102_),
    .A3(_104_),
    .B1(_109_),
    .X(_110_));
 sky130_fd_sc_hd__o32a_2 _546_ (.A1(\tcount[7] ),
    .A2(_080_),
    .A3(_085_),
    .B1(_100_),
    .B2(_110_),
    .X(sine_out[1]));
 sky130_fd_sc_hd__nand2_2 _547_ (.A(_360_),
    .B(_372_),
    .Y(_111_));
 sky130_fd_sc_hd__a21oi_2 _548_ (.A1(_037_),
    .A2(_111_),
    .B1(\tcount[3] ),
    .Y(_112_));
 sky130_fd_sc_hd__o21ai_2 _549_ (.A1(_096_),
    .A2(_112_),
    .B1(\tcount[4] ),
    .Y(_113_));
 sky130_fd_sc_hd__a21o_2 _550_ (.A1(\tcount[3] ),
    .A2(_111_),
    .B1(_105_),
    .X(_114_));
 sky130_fd_sc_hd__or3_2 _551_ (.A(\tcount[3] ),
    .B(_001_),
    .C(_353_),
    .X(_115_));
 sky130_fd_sc_hd__or2_2 _552_ (.A(_351_),
    .B(_041_),
    .X(_116_));
 sky130_fd_sc_hd__a21oi_2 _553_ (.A1(_115_),
    .A2(_116_),
    .B1(\tcount[4] ),
    .Y(_117_));
 sky130_fd_sc_hd__a41o_2 _554_ (.A1(\tcount[4] ),
    .A2(_019_),
    .A3(_041_),
    .A4(_066_),
    .B1(_117_),
    .X(_118_));
 sky130_fd_sc_hd__o211a_2 _555_ (.A1(\tcount[3] ),
    .A2(_373_),
    .B1(_063_),
    .C1(\tcount[4] ),
    .X(_119_));
 sky130_fd_sc_hd__a31o_2 _556_ (.A1(_385_),
    .A2(_039_),
    .A3(_042_),
    .B1(_348_),
    .X(_120_));
 sky130_fd_sc_hd__a221o_2 _557_ (.A1(_362_),
    .A2(_390_),
    .B1(_090_),
    .B2(_343_),
    .C1(\tcount[4] ),
    .X(_121_));
 sky130_fd_sc_hd__nand2_2 _558_ (.A(\tcount[4] ),
    .B(_361_),
    .Y(_122_));
 sky130_fd_sc_hd__o311a_2 _559_ (.A1(_344_),
    .A2(_363_),
    .A3(_122_),
    .B1(_121_),
    .C1(_031_),
    .X(_123_));
 sky130_fd_sc_hd__o221ai_2 _560_ (.A1(_052_),
    .A2(_118_),
    .B1(_119_),
    .B2(_120_),
    .C1(\tcount[7] ),
    .Y(_124_));
 sky130_fd_sc_hd__a31o_2 _561_ (.A1(_388_),
    .A2(_113_),
    .A3(_114_),
    .B1(_123_),
    .X(_125_));
 sky130_fd_sc_hd__a21oi_2 _562_ (.A1(_357_),
    .A2(_358_),
    .B1(_045_),
    .Y(_126_));
 sky130_fd_sc_hd__nor2_2 _563_ (.A(\tcount[3] ),
    .B(_072_),
    .Y(_127_));
 sky130_fd_sc_hd__and4_2 _564_ (.A(\tcount[0] ),
    .B(\tcount[3] ),
    .C(\tcount[2] ),
    .D(\tcount[1] ),
    .X(_128_));
 sky130_fd_sc_hd__or2_2 _565_ (.A(\tcount[4] ),
    .B(_128_),
    .X(_129_));
 sky130_fd_sc_hd__o221a_2 _566_ (.A1(_370_),
    .A2(_126_),
    .B1(_127_),
    .B2(_129_),
    .C1(_388_),
    .X(_130_));
 sky130_fd_sc_hd__a21oi_2 _567_ (.A1(_040_),
    .A2(_057_),
    .B1(\tcount[4] ),
    .Y(_131_));
 sky130_fd_sc_hd__a221o_2 _568_ (.A1(_022_),
    .A2(_028_),
    .B1(_040_),
    .B2(_057_),
    .C1(\tcount[4] ),
    .X(_132_));
 sky130_fd_sc_hd__or3_2 _569_ (.A(\tcount[3] ),
    .B(_045_),
    .C(_106_),
    .X(_133_));
 sky130_fd_sc_hd__and3_2 _570_ (.A(\tcount[3] ),
    .B(_356_),
    .C(_359_),
    .X(_134_));
 sky130_fd_sc_hd__or3b_2 _571_ (.A(_338_),
    .B(_349_),
    .C_N(_134_),
    .X(_135_));
 sky130_fd_sc_hd__a31o_2 _572_ (.A1(_132_),
    .A2(_133_),
    .A3(_135_),
    .B1(_348_),
    .X(_136_));
 sky130_fd_sc_hd__a221o_2 _573_ (.A1(_346_),
    .A2(_028_),
    .B1(_037_),
    .B2(\tcount[3] ),
    .C1(\tcount[4] ),
    .X(_137_));
 sky130_fd_sc_hd__or3_2 _574_ (.A(\tcount[3] ),
    .B(\tcount[1] ),
    .C(_363_),
    .X(_138_));
 sky130_fd_sc_hd__and4b_2 _575_ (.A_N(\tcount[0] ),
    .B(\tcount[3] ),
    .C(\tcount[2] ),
    .D(\tcount[1] ),
    .X(_139_));
 sky130_fd_sc_hd__or3b_2 _576_ (.A(_139_),
    .B(_338_),
    .C_N(_138_),
    .X(_140_));
 sky130_fd_sc_hd__a31o_2 _577_ (.A1(_031_),
    .A2(_137_),
    .A3(_140_),
    .B1(\tcount[7] ),
    .X(_141_));
 sky130_fd_sc_hd__or2_2 _578_ (.A(\tcount[2] ),
    .B(_041_),
    .X(_142_));
 sky130_fd_sc_hd__a211o_2 _579_ (.A1(_026_),
    .A2(_040_),
    .B1(_076_),
    .C1(\tcount[4] ),
    .X(_143_));
 sky130_fd_sc_hd__a311o_2 _580_ (.A1(_343_),
    .A2(_350_),
    .A3(_359_),
    .B1(\tcount[3] ),
    .C1(_338_),
    .X(_144_));
 sky130_fd_sc_hd__nand2_2 _581_ (.A(\tcount[4] ),
    .B(\tcount[3] ),
    .Y(_145_));
 sky130_fd_sc_hd__or3_2 _582_ (.A(_338_),
    .B(_001_),
    .C(_364_),
    .X(_146_));
 sky130_fd_sc_hd__a31o_2 _583_ (.A1(_143_),
    .A2(_144_),
    .A3(_146_),
    .B1(_052_),
    .X(_147_));
 sky130_fd_sc_hd__and4bb_2 _584_ (.A_N(_130_),
    .B_N(_141_),
    .C(_147_),
    .D(_136_),
    .X(_148_));
 sky130_fd_sc_hd__o21ba_2 _585_ (.A1(_124_),
    .A2(_125_),
    .B1_N(_148_),
    .X(sine_out[2]));
 sky130_fd_sc_hd__a211o_2 _586_ (.A1(\tcount[2] ),
    .A2(_076_),
    .B1(_126_),
    .C1(_067_),
    .X(_149_));
 sky130_fd_sc_hd__o31a_2 _587_ (.A1(\tcount[4] ),
    .A2(_363_),
    .A3(_367_),
    .B1(_149_),
    .X(_150_));
 sky130_fd_sc_hd__o211a_2 _588_ (.A1(_364_),
    .A2(_373_),
    .B1(_092_),
    .C1(\tcount[4] ),
    .X(_151_));
 sky130_fd_sc_hd__nand2_2 _589_ (.A(_345_),
    .B(_028_),
    .Y(_152_));
 sky130_fd_sc_hd__a31o_2 _590_ (.A1(_338_),
    .A2(_037_),
    .A3(_152_),
    .B1(_348_),
    .X(_153_));
 sky130_fd_sc_hd__a32o_2 _591_ (.A1(\tcount[3] ),
    .A2(\tcount[1] ),
    .A3(_026_),
    .B1(_076_),
    .B2(_360_),
    .X(_154_));
 sky130_fd_sc_hd__nand2_2 _592_ (.A(\tcount[4] ),
    .B(_154_),
    .Y(_155_));
 sky130_fd_sc_hd__a21oi_2 _593_ (.A1(\tcount[0] ),
    .A2(\tcount[2] ),
    .B1(\tcount[3] ),
    .Y(_156_));
 sky130_fd_sc_hd__nand2_2 _594_ (.A(_346_),
    .B(_156_),
    .Y(_157_));
 sky130_fd_sc_hd__a31o_2 _595_ (.A1(_023_),
    .A2(_063_),
    .A3(_157_),
    .B1(\tcount[4] ),
    .X(_158_));
 sky130_fd_sc_hd__a21o_2 _596_ (.A1(_155_),
    .A2(_158_),
    .B1(_389_),
    .X(_159_));
 sky130_fd_sc_hd__o31a_2 _597_ (.A1(_339_),
    .A2(_045_),
    .A3(_056_),
    .B1(_083_),
    .X(_160_));
 sky130_fd_sc_hd__a21oi_2 _598_ (.A1(_368_),
    .A2(_037_),
    .B1(_339_),
    .Y(_161_));
 sky130_fd_sc_hd__a211o_2 _599_ (.A1(\tcount[2] ),
    .A2(_076_),
    .B1(_161_),
    .C1(_067_),
    .X(_162_));
 sky130_fd_sc_hd__a21oi_2 _600_ (.A1(\tcount[4] ),
    .A2(_162_),
    .B1(_160_),
    .Y(_163_));
 sky130_fd_sc_hd__o21a_2 _601_ (.A1(_052_),
    .A2(_150_),
    .B1(_159_),
    .X(_164_));
 sky130_fd_sc_hd__o221a_2 _602_ (.A1(_151_),
    .A2(_153_),
    .B1(_163_),
    .B2(_032_),
    .C1(\tcount[7] ),
    .X(_165_));
 sky130_fd_sc_hd__or2_2 _603_ (.A(_344_),
    .B(_082_),
    .X(_166_));
 sky130_fd_sc_hd__a311o_2 _604_ (.A1(\tcount[4] ),
    .A2(_042_),
    .A3(_166_),
    .B1(_160_),
    .C1(_032_),
    .X(_167_));
 sky130_fd_sc_hd__or2_2 _605_ (.A(\tcount[4] ),
    .B(_072_),
    .X(_168_));
 sky130_fd_sc_hd__a31o_2 _606_ (.A1(_051_),
    .A2(_149_),
    .A3(_168_),
    .B1(\tcount[7] ),
    .X(_169_));
 sky130_fd_sc_hd__o31a_2 _607_ (.A1(_339_),
    .A2(_367_),
    .A3(_025_),
    .B1(_092_),
    .X(_170_));
 sky130_fd_sc_hd__a221o_2 _608_ (.A1(\tcount[3] ),
    .A2(_037_),
    .B1(_057_),
    .B2(_372_),
    .C1(\tcount[4] ),
    .X(_171_));
 sky130_fd_sc_hd__o211a_2 _609_ (.A1(_338_),
    .A2(_170_),
    .B1(_171_),
    .C1(_347_),
    .X(_172_));
 sky130_fd_sc_hd__o21a_2 _610_ (.A1(_000_),
    .A2(_376_),
    .B1(_065_),
    .X(_173_));
 sky130_fd_sc_hd__o211a_2 _611_ (.A1(\tcount[4] ),
    .A2(_173_),
    .B1(_155_),
    .C1(_388_),
    .X(_174_));
 sky130_fd_sc_hd__or3b_2 _612_ (.A(_169_),
    .B(_172_),
    .C_N(_167_),
    .X(_175_));
 sky130_fd_sc_hd__o2bb2a_2 _613_ (.A1_N(_164_),
    .A2_N(_165_),
    .B1(_174_),
    .B2(_175_),
    .X(sine_out[3]));
 sky130_fd_sc_hd__nor2_2 _614_ (.A(_027_),
    .B(_107_),
    .Y(_176_));
 sky130_fd_sc_hd__or3b_2 _615_ (.A(_339_),
    .B(_360_),
    .C_N(_386_),
    .X(_177_));
 sky130_fd_sc_hd__o211a_2 _616_ (.A1(_338_),
    .A2(_176_),
    .B1(_177_),
    .C1(_388_),
    .X(_178_));
 sky130_fd_sc_hd__nand2_2 _617_ (.A(_345_),
    .B(_064_),
    .Y(_179_));
 sky130_fd_sc_hd__o21a_2 _618_ (.A1(\tcount[2] ),
    .A2(_346_),
    .B1(_156_),
    .X(_180_));
 sky130_fd_sc_hd__a31o_2 _619_ (.A1(\tcount[0] ),
    .A2(\tcount[3] ),
    .A3(\tcount[2] ),
    .B1(\tcount[4] ),
    .X(_181_));
 sky130_fd_sc_hd__o32ai_2 _620_ (.A1(_338_),
    .A2(_060_),
    .A3(_161_),
    .B1(_180_),
    .B2(_181_),
    .Y(_182_));
 sky130_fd_sc_hd__nor2_2 _621_ (.A(_379_),
    .B(_064_),
    .Y(_183_));
 sky130_fd_sc_hd__a31o_2 _622_ (.A1(_338_),
    .A2(_377_),
    .A3(_183_),
    .B1(\tcount[5] ),
    .X(_184_));
 sky130_fd_sc_hd__nor4_2 _623_ (.A(_338_),
    .B(_380_),
    .C(_082_),
    .D(_139_),
    .Y(_185_));
 sky130_fd_sc_hd__a311o_2 _624_ (.A1(_338_),
    .A2(_377_),
    .A3(_183_),
    .B1(_185_),
    .C1(\tcount[5] ),
    .X(_186_));
 sky130_fd_sc_hd__a21bo_2 _625_ (.A1(\tcount[2] ),
    .A2(_076_),
    .B1_N(_364_),
    .X(_187_));
 sky130_fd_sc_hd__a221o_2 _626_ (.A1(_029_),
    .A2(_049_),
    .B1(_187_),
    .B2(\tcount[4] ),
    .C1(_337_),
    .X(_188_));
 sky130_fd_sc_hd__a32o_2 _627_ (.A1(\tcount[6] ),
    .A2(_186_),
    .A3(_188_),
    .B1(_051_),
    .B2(_182_),
    .X(_189_));
 sky130_fd_sc_hd__a21oi_2 _628_ (.A1(_178_),
    .A2(_179_),
    .B1(_189_),
    .Y(_190_));
 sky130_fd_sc_hd__or3_2 _629_ (.A(\tcount[7] ),
    .B(_178_),
    .C(_189_),
    .X(_191_));
 sky130_fd_sc_hd__o21ai_2 _630_ (.A1(_341_),
    .A2(_190_),
    .B1(_191_),
    .Y(sine_out[4]));
 sky130_fd_sc_hd__o22a_2 _631_ (.A1(\tcount[0] ),
    .A2(_360_),
    .B1(_361_),
    .B2(_089_),
    .X(_192_));
 sky130_fd_sc_hd__o21ai_2 _632_ (.A1(_044_),
    .A2(_192_),
    .B1(\tcount[4] ),
    .Y(_193_));
 sky130_fd_sc_hd__a31o_2 _633_ (.A1(\tcount[3] ),
    .A2(_343_),
    .A3(_037_),
    .B1(\tcount[4] ),
    .X(_194_));
 sky130_fd_sc_hd__or2_2 _634_ (.A(_047_),
    .B(_194_),
    .X(_195_));
 sky130_fd_sc_hd__a21oi_2 _635_ (.A1(_193_),
    .A2(_195_),
    .B1(_389_),
    .Y(_196_));
 sky130_fd_sc_hd__o211a_2 _636_ (.A1(\tcount[0] ),
    .A2(_360_),
    .B1(_022_),
    .C1(_356_),
    .X(_197_));
 sky130_fd_sc_hd__a221o_2 _637_ (.A1(\tcount[0] ),
    .A2(_354_),
    .B1(_359_),
    .B2(_069_),
    .C1(\tcount[3] ),
    .X(_198_));
 sky130_fd_sc_hd__a311o_2 _638_ (.A1(_354_),
    .A2(_356_),
    .A3(_198_),
    .B1(_067_),
    .C1(_338_),
    .X(_199_));
 sky130_fd_sc_hd__o311a_2 _639_ (.A1(\tcount[4] ),
    .A2(_048_),
    .A3(_058_),
    .B1(_199_),
    .C1(_031_),
    .X(_200_));
 sky130_fd_sc_hd__o311a_2 _640_ (.A1(\tcount[3] ),
    .A2(_353_),
    .A3(_025_),
    .B1(_361_),
    .C1(\tcount[4] ),
    .X(_201_));
 sky130_fd_sc_hd__or3_2 _641_ (.A(_339_),
    .B(_351_),
    .C(_036_),
    .X(_202_));
 sky130_fd_sc_hd__a21oi_2 _642_ (.A1(_115_),
    .A2(_202_),
    .B1(\tcount[4] ),
    .Y(_203_));
 sky130_fd_sc_hd__o21a_2 _643_ (.A1(_201_),
    .A2(_203_),
    .B1(_347_),
    .X(_204_));
 sky130_fd_sc_hd__o21a_2 _644_ (.A1(_355_),
    .A2(_361_),
    .B1(_338_),
    .X(_205_));
 sky130_fd_sc_hd__a32o_2 _645_ (.A1(\tcount[4] ),
    .A2(_063_),
    .A3(_198_),
    .B1(_205_),
    .B2(_369_),
    .X(_206_));
 sky130_fd_sc_hd__nand2_2 _646_ (.A(_051_),
    .B(_206_),
    .Y(_207_));
 sky130_fd_sc_hd__or4b_2 _647_ (.A(_196_),
    .B(_200_),
    .C(_204_),
    .D_N(_207_),
    .X(_208_));
 sky130_fd_sc_hd__a21o_2 _648_ (.A1(\tcount[0] ),
    .A2(_018_),
    .B1(_194_),
    .X(_209_));
 sky130_fd_sc_hd__a21o_2 _649_ (.A1(_193_),
    .A2(_209_),
    .B1(_389_),
    .X(_210_));
 sky130_fd_sc_hd__and4bb_2 _650_ (.A_N(_200_),
    .B_N(_204_),
    .C(_207_),
    .D(_210_),
    .X(_211_));
 sky130_fd_sc_hd__mux2_1 _651_ (.A0(_208_),
    .A1(_211_),
    .S(_341_),
    .X(sine_out[5]));
 sky130_fd_sc_hd__a21oi_2 _652_ (.A1(\tcount[1] ),
    .A2(_156_),
    .B1(_103_),
    .Y(_212_));
 sky130_fd_sc_hd__o21a_2 _653_ (.A1(_087_),
    .A2(_112_),
    .B1(_338_),
    .X(_213_));
 sky130_fd_sc_hd__o21ai_2 _654_ (.A1(_212_),
    .A2(_213_),
    .B1(_388_),
    .Y(_214_));
 sky130_fd_sc_hd__o211a_2 _655_ (.A1(\tcount[3] ),
    .A2(_366_),
    .B1(_377_),
    .C1(\tcount[4] ),
    .X(_215_));
 sky130_fd_sc_hd__nand2_2 _656_ (.A(_037_),
    .B(_076_),
    .Y(_216_));
 sky130_fd_sc_hd__and3_2 _657_ (.A(_338_),
    .B(_202_),
    .C(_216_),
    .X(_217_));
 sky130_fd_sc_hd__or3_2 _658_ (.A(_032_),
    .B(_215_),
    .C(_217_),
    .X(_218_));
 sky130_fd_sc_hd__a32o_2 _659_ (.A1(\tcount[3] ),
    .A2(_352_),
    .A3(_022_),
    .B1(_358_),
    .B2(_340_),
    .X(_219_));
 sky130_fd_sc_hd__a22o_2 _660_ (.A1(_029_),
    .A2(_042_),
    .B1(_219_),
    .B2(\tcount[4] ),
    .X(_220_));
 sky130_fd_sc_hd__a211o_2 _661_ (.A1(\tcount[2] ),
    .A2(_001_),
    .B1(_036_),
    .C1(_339_),
    .X(_221_));
 sky130_fd_sc_hd__a22o_2 _662_ (.A1(\tcount[3] ),
    .A2(_372_),
    .B1(_037_),
    .B2(_076_),
    .X(_222_));
 sky130_fd_sc_hd__a22o_2 _663_ (.A1(_083_),
    .A2(_221_),
    .B1(_222_),
    .B2(\tcount[4] ),
    .X(_223_));
 sky130_fd_sc_hd__o2bb2a_2 _664_ (.A1_N(_051_),
    .A2_N(_220_),
    .B1(_223_),
    .B2(_348_),
    .X(_224_));
 sky130_fd_sc_hd__and3_2 _665_ (.A(\tcount[7] ),
    .B(_218_),
    .C(_224_),
    .X(_225_));
 sky130_fd_sc_hd__o21ai_2 _666_ (.A1(_215_),
    .A2(_217_),
    .B1(_031_),
    .Y(_226_));
 sky130_fd_sc_hd__nand2_2 _667_ (.A(_347_),
    .B(_223_),
    .Y(_227_));
 sky130_fd_sc_hd__a311o_2 _668_ (.A1(_338_),
    .A2(_381_),
    .A3(_142_),
    .B1(_212_),
    .C1(_389_),
    .X(_228_));
 sky130_fd_sc_hd__o2111a_2 _669_ (.A1(_052_),
    .A2(_220_),
    .B1(_226_),
    .C1(_227_),
    .D1(_228_),
    .X(_229_));
 sky130_fd_sc_hd__a22oi_2 _670_ (.A1(_214_),
    .A2(_225_),
    .B1(_229_),
    .B2(_341_),
    .Y(sine_out[6]));
 sky130_fd_sc_hd__or2_2 _671_ (.A(_344_),
    .B(_364_),
    .X(_230_));
 sky130_fd_sc_hd__nand2_2 _672_ (.A(\tcount[4] ),
    .B(_066_),
    .Y(_231_));
 sky130_fd_sc_hd__a2bb2o_2 _673_ (.A1_N(_366_),
    .A2_N(_231_),
    .B1(_230_),
    .B2(_385_),
    .X(_232_));
 sky130_fd_sc_hd__a221o_2 _674_ (.A1(_339_),
    .A2(_072_),
    .B1(_074_),
    .B2(_354_),
    .C1(\tcount[4] ),
    .X(_233_));
 sky130_fd_sc_hd__nor2_2 _675_ (.A(\tcount[2] ),
    .B(_039_),
    .Y(_234_));
 sky130_fd_sc_hd__a211o_2 _676_ (.A1(_345_),
    .A2(_107_),
    .B1(_234_),
    .C1(_338_),
    .X(_235_));
 sky130_fd_sc_hd__a32o_2 _677_ (.A1(_031_),
    .A2(_233_),
    .A3(_235_),
    .B1(_232_),
    .B2(_347_),
    .X(_236_));
 sky130_fd_sc_hd__or3_2 _678_ (.A(_338_),
    .B(_379_),
    .C(_380_),
    .X(_237_));
 sky130_fd_sc_hd__a31o_2 _679_ (.A1(\tcount[3] ),
    .A2(_027_),
    .A3(_072_),
    .B1(_237_),
    .X(_238_));
 sky130_fd_sc_hd__a311o_2 _680_ (.A1(\tcount[3] ),
    .A2(_354_),
    .A3(_356_),
    .B1(_046_),
    .C1(\tcount[4] ),
    .X(_239_));
 sky130_fd_sc_hd__a31o_2 _681_ (.A1(_331_),
    .A2(_238_),
    .A3(_239_),
    .B1(_388_),
    .X(_240_));
 sky130_fd_sc_hd__o21a_2 _682_ (.A1(_045_),
    .A2(_069_),
    .B1(\tcount[3] ),
    .X(_241_));
 sky130_fd_sc_hd__o21ai_2 _683_ (.A1(_059_),
    .A2(_241_),
    .B1(\tcount[4] ),
    .Y(_242_));
 sky130_fd_sc_hd__or4_2 _684_ (.A(\tcount[4] ),
    .B(_349_),
    .C(_363_),
    .D(_384_),
    .X(_243_));
 sky130_fd_sc_hd__a21o_2 _685_ (.A1(_242_),
    .A2(_243_),
    .B1(\tcount[5] ),
    .X(_244_));
 sky130_fd_sc_hd__nand2_2 _686_ (.A(_385_),
    .B(_142_),
    .Y(_245_));
 sky130_fd_sc_hd__a21o_2 _687_ (.A1(_242_),
    .A2(_245_),
    .B1(\tcount[5] ),
    .X(_246_));
 sky130_fd_sc_hd__a21oi_2 _688_ (.A1(_240_),
    .A2(_246_),
    .B1(_236_),
    .Y(_247_));
 sky130_fd_sc_hd__a211o_2 _689_ (.A1(_240_),
    .A2(_244_),
    .B1(_341_),
    .C1(_236_),
    .X(_248_));
 sky130_fd_sc_hd__o21ai_2 _690_ (.A1(\tcount[7] ),
    .A2(_247_),
    .B1(_248_),
    .Y(sine_out[7]));
 sky130_fd_sc_hd__or3_2 _691_ (.A(_338_),
    .B(\tcount[3] ),
    .C(_070_),
    .X(_249_));
 sky130_fd_sc_hd__o41a_2 _692_ (.A1(_338_),
    .A2(\tcount[1] ),
    .A3(_363_),
    .A4(_018_),
    .B1(_249_),
    .X(_250_));
 sky130_fd_sc_hd__and3_2 _693_ (.A(\tcount[3] ),
    .B(_345_),
    .C(_026_),
    .X(_251_));
 sky130_fd_sc_hd__o31ai_2 _694_ (.A1(\tcount[4] ),
    .A2(_047_),
    .A3(_251_),
    .B1(_250_),
    .Y(_252_));
 sky130_fd_sc_hd__or3_2 _695_ (.A(_338_),
    .B(_047_),
    .C(_241_),
    .X(_253_));
 sky130_fd_sc_hd__a21o_2 _696_ (.A1(_339_),
    .A2(_390_),
    .B1(\tcount[4] ),
    .X(_254_));
 sky130_fd_sc_hd__a21o_2 _697_ (.A1(\tcount[3] ),
    .A2(_197_),
    .B1(_254_),
    .X(_255_));
 sky130_fd_sc_hd__a31o_2 _698_ (.A1(_340_),
    .A2(_066_),
    .A3(_107_),
    .B1(\tcount[4] ),
    .X(_256_));
 sky130_fd_sc_hd__or3_2 _699_ (.A(_339_),
    .B(_355_),
    .C(_106_),
    .X(_257_));
 sky130_fd_sc_hd__a31oi_2 _700_ (.A1(_249_),
    .A2(_256_),
    .A3(_257_),
    .B1(_052_),
    .Y(_258_));
 sky130_fd_sc_hd__a21oi_2 _701_ (.A1(_346_),
    .A2(_065_),
    .B1(_371_),
    .Y(_259_));
 sky130_fd_sc_hd__and3b_2 _702_ (.A_N(\tcount[2] ),
    .B(\tcount[3] ),
    .C(\tcount[0] ),
    .X(_260_));
 sky130_fd_sc_hd__o21ai_2 _703_ (.A1(_342_),
    .A2(_026_),
    .B1(\tcount[3] ),
    .Y(_261_));
 sky130_fd_sc_hd__a311o_2 _704_ (.A1(\tcount[3] ),
    .A2(_354_),
    .A3(_356_),
    .B1(_260_),
    .C1(\tcount[4] ),
    .X(_262_));
 sky130_fd_sc_hd__o311a_2 _705_ (.A1(_338_),
    .A2(_074_),
    .A3(_259_),
    .B1(_262_),
    .C1(_347_),
    .X(_263_));
 sky130_fd_sc_hd__a31o_2 _706_ (.A1(_031_),
    .A2(_253_),
    .A3(_255_),
    .B1(_263_),
    .X(_264_));
 sky130_fd_sc_hd__a211o_2 _707_ (.A1(_388_),
    .A2(_252_),
    .B1(_258_),
    .C1(_264_),
    .X(_265_));
 sky130_fd_sc_hd__a211o_2 _708_ (.A1(\tcount[0] ),
    .A2(_018_),
    .B1(_251_),
    .C1(\tcount[4] ),
    .X(_266_));
 sky130_fd_sc_hd__a21oi_2 _709_ (.A1(_250_),
    .A2(_266_),
    .B1(_389_),
    .Y(_267_));
 sky130_fd_sc_hd__or4_2 _710_ (.A(\tcount[7] ),
    .B(_258_),
    .C(_264_),
    .D(_267_),
    .X(_268_));
 sky130_fd_sc_hd__a21bo_2 _711_ (.A1(\tcount[7] ),
    .A2(_265_),
    .B1_N(_268_),
    .X(sine_out[8]));
 sky130_fd_sc_hd__nand2_2 _712_ (.A(_001_),
    .B(_018_),
    .Y(_269_));
 sky130_fd_sc_hd__a21o_2 _713_ (.A1(_261_),
    .A2(_269_),
    .B1(_338_),
    .X(_270_));
 sky130_fd_sc_hd__o31a_2 _714_ (.A1(\tcount[4] ),
    .A2(_020_),
    .A3(_096_),
    .B1(_270_),
    .X(_271_));
 sky130_fd_sc_hd__a31o_2 _715_ (.A1(\tcount[4] ),
    .A2(_071_),
    .A3(_198_),
    .B1(_348_),
    .X(_272_));
 sky130_fd_sc_hd__o221a_2 _716_ (.A1(_355_),
    .A2(_364_),
    .B1(_069_),
    .B2(\tcount[3] ),
    .C1(_338_),
    .X(_273_));
 sky130_fd_sc_hd__a311o_2 _717_ (.A1(\tcount[4] ),
    .A2(_138_),
    .A3(_142_),
    .B1(_273_),
    .C1(_052_),
    .X(_274_));
 sky130_fd_sc_hd__nand2_2 _718_ (.A(\tcount[3] ),
    .B(_346_),
    .Y(_275_));
 sky130_fd_sc_hd__o221a_2 _719_ (.A1(_361_),
    .A2(_367_),
    .B1(_019_),
    .B2(_346_),
    .C1(\tcount[4] ),
    .X(_276_));
 sky130_fd_sc_hd__a311o_2 _720_ (.A1(_338_),
    .A2(_025_),
    .A3(_275_),
    .B1(_276_),
    .C1(_032_),
    .X(_277_));
 sky130_fd_sc_hd__o211a_2 _721_ (.A1(_131_),
    .A2(_272_),
    .B1(_274_),
    .C1(_277_),
    .X(_278_));
 sky130_fd_sc_hd__a211o_2 _722_ (.A1(_018_),
    .A2(_057_),
    .B1(_096_),
    .C1(\tcount[4] ),
    .X(_279_));
 sky130_fd_sc_hd__a21o_2 _723_ (.A1(_270_),
    .A2(_279_),
    .B1(_389_),
    .X(_280_));
 sky130_fd_sc_hd__nand2_2 _724_ (.A(_278_),
    .B(_280_),
    .Y(_281_));
 sky130_fd_sc_hd__o211a_2 _725_ (.A1(_389_),
    .A2(_271_),
    .B1(_278_),
    .C1(_341_),
    .X(_282_));
 sky130_fd_sc_hd__a21o_2 _726_ (.A1(\tcount[7] ),
    .A2(_281_),
    .B1(_282_),
    .X(sine_out[9]));
 sky130_fd_sc_hd__o41a_2 _727_ (.A1(\tcount[3] ),
    .A2(_342_),
    .A3(_351_),
    .A4(_367_),
    .B1(_357_),
    .X(_283_));
 sky130_fd_sc_hd__a21o_2 _728_ (.A1(_343_),
    .A2(_374_),
    .B1(\tcount[4] ),
    .X(_284_));
 sky130_fd_sc_hd__o211ai_2 _729_ (.A1(_338_),
    .A2(_283_),
    .B1(_284_),
    .C1(_347_),
    .Y(_285_));
 sky130_fd_sc_hd__o221a_2 _730_ (.A1(_373_),
    .A2(_019_),
    .B1(_075_),
    .B2(_353_),
    .C1(_338_),
    .X(_286_));
 sky130_fd_sc_hd__a211o_2 _731_ (.A1(\tcount[2] ),
    .A2(_001_),
    .B1(_349_),
    .C1(_371_),
    .X(_287_));
 sky130_fd_sc_hd__o211a_2 _732_ (.A1(\tcount[3] ),
    .A2(_197_),
    .B1(_287_),
    .C1(\tcount[4] ),
    .X(_288_));
 sky130_fd_sc_hd__o31a_2 _733_ (.A1(_032_),
    .A2(_286_),
    .A3(_288_),
    .B1(_285_),
    .X(_289_));
 sky130_fd_sc_hd__nand2_2 _734_ (.A(_372_),
    .B(_028_),
    .Y(_290_));
 sky130_fd_sc_hd__a21oi_2 _735_ (.A1(_001_),
    .A2(_023_),
    .B1(_129_),
    .Y(_291_));
 sky130_fd_sc_hd__a211o_2 _736_ (.A1(\tcount[4] ),
    .A2(_290_),
    .B1(_291_),
    .C1(_052_),
    .X(_292_));
 sky130_fd_sc_hd__nand2_2 _737_ (.A(_372_),
    .B(_076_),
    .Y(_293_));
 sky130_fd_sc_hd__or2_2 _738_ (.A(_338_),
    .B(_384_),
    .X(_294_));
 sky130_fd_sc_hd__a31o_2 _739_ (.A1(_037_),
    .A2(_111_),
    .A3(_293_),
    .B1(_294_),
    .X(_295_));
 sky130_fd_sc_hd__or4_2 _740_ (.A(\tcount[4] ),
    .B(_351_),
    .C(_384_),
    .D(_260_),
    .X(_296_));
 sky130_fd_sc_hd__a21o_2 _741_ (.A1(_295_),
    .A2(_296_),
    .B1(_389_),
    .X(_297_));
 sky130_fd_sc_hd__and3_2 _742_ (.A(_289_),
    .B(_292_),
    .C(_297_),
    .X(_298_));
 sky130_fd_sc_hd__or3_2 _743_ (.A(\tcount[4] ),
    .B(_069_),
    .C(_092_),
    .X(_299_));
 sky130_fd_sc_hd__or3_2 _744_ (.A(\tcount[4] ),
    .B(_339_),
    .C(_026_),
    .X(_300_));
 sky130_fd_sc_hd__a31o_2 _745_ (.A1(_295_),
    .A2(_299_),
    .A3(_300_),
    .B1(_389_),
    .X(_301_));
 sky130_fd_sc_hd__and3_2 _746_ (.A(\tcount[7] ),
    .B(_289_),
    .C(_292_),
    .X(_302_));
 sky130_fd_sc_hd__o2bb2a_2 _747_ (.A1_N(_301_),
    .A2_N(_302_),
    .B1(\tcount[7] ),
    .B2(_298_),
    .X(sine_out[10]));
 sky130_fd_sc_hd__or3b_2 _748_ (.A(_161_),
    .B(_294_),
    .C_N(_179_),
    .X(_303_));
 sky130_fd_sc_hd__a31o_2 _749_ (.A1(_016_),
    .A2(_023_),
    .A3(_063_),
    .B1(\tcount[4] ),
    .X(_304_));
 sky130_fd_sc_hd__o2111a_2 _750_ (.A1(_374_),
    .A2(_090_),
    .B1(_035_),
    .C1(_337_),
    .D1(\tcount[4] ),
    .X(_305_));
 sky130_fd_sc_hd__a311o_2 _751_ (.A1(\tcount[5] ),
    .A2(_303_),
    .A3(_304_),
    .B1(_305_),
    .C1(_331_),
    .X(_306_));
 sky130_fd_sc_hd__a211o_2 _752_ (.A1(_360_),
    .A2(_372_),
    .B1(_082_),
    .C1(\tcount[4] ),
    .X(_307_));
 sky130_fd_sc_hd__nand2_2 _753_ (.A(\tcount[4] ),
    .B(_065_),
    .Y(_308_));
 sky130_fd_sc_hd__a31oi_2 _754_ (.A1(\tcount[5] ),
    .A2(_307_),
    .A3(_308_),
    .B1(\tcount[6] ),
    .Y(_309_));
 sky130_fd_sc_hd__a21o_2 _755_ (.A1(_368_),
    .A2(_037_),
    .B1(\tcount[3] ),
    .X(_310_));
 sky130_fd_sc_hd__o311a_2 _756_ (.A1(_339_),
    .A2(_367_),
    .A3(_036_),
    .B1(_086_),
    .C1(\tcount[4] ),
    .X(_311_));
 sky130_fd_sc_hd__a311o_2 _757_ (.A1(_338_),
    .A2(_377_),
    .A3(_310_),
    .B1(_311_),
    .C1(\tcount[5] ),
    .X(_312_));
 sky130_fd_sc_hd__nand2_2 _758_ (.A(_309_),
    .B(_312_),
    .Y(_313_));
 sky130_fd_sc_hd__o21ai_2 _759_ (.A1(_184_),
    .A2(_311_),
    .B1(_309_),
    .Y(_314_));
 sky130_fd_sc_hd__a21oi_2 _760_ (.A1(_306_),
    .A2(_314_),
    .B1(\tcount[7] ),
    .Y(_315_));
 sky130_fd_sc_hd__a31o_2 _761_ (.A1(\tcount[7] ),
    .A2(_306_),
    .A3(_313_),
    .B1(_315_),
    .X(sine_out[11]));
 sky130_fd_sc_hd__a211o_2 _762_ (.A1(\tcount[0] ),
    .A2(_384_),
    .B1(_134_),
    .C1(\tcount[4] ),
    .X(_316_));
 sky130_fd_sc_hd__o31ai_2 _763_ (.A1(_349_),
    .A2(_363_),
    .A3(_134_),
    .B1(\tcount[4] ),
    .Y(_317_));
 sky130_fd_sc_hd__a31o_2 _764_ (.A1(_337_),
    .A2(\tcount[4] ),
    .A3(_091_),
    .B1(_331_),
    .X(_318_));
 sky130_fd_sc_hd__a31o_2 _765_ (.A1(\tcount[5] ),
    .A2(_316_),
    .A3(_317_),
    .B1(_318_),
    .X(_319_));
 sky130_fd_sc_hd__a22o_2 _766_ (.A1(\tcount[3] ),
    .A2(_359_),
    .B1(_076_),
    .B2(\tcount[2] ),
    .X(_320_));
 sky130_fd_sc_hd__and2_2 _767_ (.A(_338_),
    .B(_320_),
    .X(_321_));
 sky130_fd_sc_hd__a21oi_2 _768_ (.A1(\tcount[4] ),
    .A2(_350_),
    .B1(_134_),
    .Y(_322_));
 sky130_fd_sc_hd__a31o_2 _769_ (.A1(\tcount[4] ),
    .A2(\tcount[3] ),
    .A3(_359_),
    .B1(_389_),
    .X(_323_));
 sky130_fd_sc_hd__o221a_2 _770_ (.A1(_052_),
    .A2(_321_),
    .B1(_322_),
    .B2(_323_),
    .C1(_319_),
    .X(_324_));
 sky130_fd_sc_hd__or2_2 _771_ (.A(\tcount[4] ),
    .B(_179_),
    .X(_325_));
 sky130_fd_sc_hd__and2_2 _772_ (.A(\tcount[7] ),
    .B(_325_),
    .X(_326_));
 sky130_fd_sc_hd__mux2_1 _773_ (.A0(_341_),
    .A1(_326_),
    .S(_324_),
    .X(sine_out[12]));
 sky130_fd_sc_hd__a22o_2 _774_ (.A1(_051_),
    .A2(_183_),
    .B1(_284_),
    .B2(_145_),
    .X(_327_));
 sky130_fd_sc_hd__or2_2 _775_ (.A(_347_),
    .B(_327_),
    .X(_328_));
 sky130_fd_sc_hd__o21a_2 _776_ (.A1(\tcount[5] ),
    .A2(_325_),
    .B1(\tcount[7] ),
    .X(_329_));
 sky130_fd_sc_hd__mux2_1 _777_ (.A0(_329_),
    .A1(_341_),
    .S(_328_),
    .X(sine_out[13]));
 sky130_fd_sc_hd__a32oi_2 _778_ (.A1(_388_),
    .A2(_145_),
    .A3(_325_),
    .B1(_284_),
    .B2(_031_),
    .Y(_330_));
 sky130_fd_sc_hd__or3_2 _779_ (.A(\tcount[6] ),
    .B(\tcount[5] ),
    .C(_325_),
    .X(_332_));
 sky130_fd_sc_hd__a21oi_2 _780_ (.A1(_330_),
    .A2(_332_),
    .B1(\tcount[7] ),
    .Y(_333_));
 sky130_fd_sc_hd__a21oi_2 _781_ (.A1(\tcount[7] ),
    .A2(_330_),
    .B1(_333_),
    .Y(sine_out[14]));
 sky130_fd_sc_hd__and2_2 _782_ (.A(\tcount[7] ),
    .B(_332_),
    .X(sine_out[15]));
 sky130_fd_sc_hd__nor2_2 _783_ (.A(_090_),
    .B(_128_),
    .Y(_003_));
 sky130_fd_sc_hd__nand2_2 _784_ (.A(\tcount[4] ),
    .B(_128_),
    .Y(_334_));
 sky130_fd_sc_hd__and2_2 _785_ (.A(_129_),
    .B(_334_),
    .X(_004_));
 sky130_fd_sc_hd__xnor2_2 _786_ (.A(\tcount[5] ),
    .B(_334_),
    .Y(_005_));
 sky130_fd_sc_hd__or2_2 _787_ (.A(_032_),
    .B(_334_),
    .X(_335_));
 sky130_fd_sc_hd__a31o_2 _788_ (.A1(\tcount[5] ),
    .A2(\tcount[4] ),
    .A3(_128_),
    .B1(\tcount[6] ),
    .X(_336_));
 sky130_fd_sc_hd__and2_2 _789_ (.A(_335_),
    .B(_336_),
    .X(_006_));
 sky130_fd_sc_hd__xnor2_2 _790_ (.A(\tcount[7] ),
    .B(_335_),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _791_ (.A(rst),
    .Y(_009_));
 sky130_fd_sc_hd__inv_2 _792_ (.A(rst),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _793_ (.A(rst),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _794_ (.A(rst),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _795_ (.A(rst),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _796_ (.A(rst),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _797_ (.A(rst),
    .Y(_015_));
 sky130_fd_sc_hd__dfrtp_2 _798_ (.CLK(clk),
    .D(_000_),
    .RESET_B(_008_),
    .Q(\tcount[0] ));
 sky130_fd_sc_hd__dfrtp_2 _799_ (.CLK(clk),
    .D(_001_),
    .RESET_B(_009_),
    .Q(\tcount[1] ));
 sky130_fd_sc_hd__dfrtp_2 _800_ (.CLK(clk),
    .D(_002_),
    .RESET_B(_010_),
    .Q(\tcount[2] ));
 sky130_fd_sc_hd__dfrtp_2 _801_ (.CLK(clk),
    .D(_003_),
    .RESET_B(_011_),
    .Q(\tcount[3] ));
 sky130_fd_sc_hd__dfrtp_2 _802_ (.CLK(clk),
    .D(_004_),
    .RESET_B(_012_),
    .Q(\tcount[4] ));
 sky130_fd_sc_hd__dfrtp_2 _803_ (.CLK(clk),
    .D(_005_),
    .RESET_B(_013_),
    .Q(\tcount[5] ));
 sky130_fd_sc_hd__dfrtp_2 _804_ (.CLK(clk),
    .D(_006_),
    .RESET_B(_014_),
    .Q(\tcount[6] ));
 sky130_fd_sc_hd__dfrtp_2 _805_ (.CLK(clk),
    .D(_007_),
    .RESET_B(_015_),
    .Q(\tcount[7] ));
endmodule
