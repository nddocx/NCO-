* NGSPICE file created from counter_8bit.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

.subckt counter_8bit VGND VPWR clk rst sine_out[0] sine_out[10] sine_out[11] sine_out[12]
+ sine_out[13] sine_out[14] sine_out[15] sine_out[1] sine_out[2] sine_out[3] sine_out[4]
+ sine_out[5] sine_out[6] sine_out[7] sine_out[8] sine_out[9]
XTAP_TAPCELL_ROW_24_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_432_ net47 net58 VGND VGND VPWR VPWR _374_ sky130_fd_sc_hd__and2_1
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_501_ net46 net67 VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__nand2b_1
XFILLER_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_415_ net65 net51 VGND VGND VPWR VPWR _357_ sky130_fd_sc_hd__nand2b_1
XFILLER_23_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_680_ net48 _354_ _356_ _046_ net41 VGND VGND VPWR VPWR _239_ sky130_fd_sc_hd__a311o_1
XFILLER_29_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_801_ clknet_1_0__leaf_clk _003_ _011_ VGND VGND VPWR VPWR tcount\[3\] sky130_fd_sc_hd__dfrtp_1
X_594_ net23 _156_ VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__nand2_1
X_663_ _083_ _221_ _222_ net38 VGND VGND VPWR VPWR _223_ sky130_fd_sc_hd__a22o_1
X_732_ net45 _197_ _287_ net35 VGND VGND VPWR VPWR _288_ sky130_fd_sc_hd__o211a_1
XFILLER_19_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput7 net7 VGND VGND VPWR VPWR sine_out[14] sky130_fd_sc_hd__buf_2
X_646_ _051_ _206_ VGND VGND VPWR VPWR _207_ sky130_fd_sc_hd__nand2_1
XFILLER_16_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_577_ _031_ _137_ _140_ net31 VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__a31o_1
X_715_ net36 _071_ _198_ _348_ VGND VGND VPWR VPWR _272_ sky130_fd_sc_hd__a31o_1
X_500_ net52 net61 VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__or2_2
X_431_ net59 net23 VGND VGND VPWR VPWR _373_ sky130_fd_sc_hd__and2_1
X_629_ net31 _178_ _189_ VGND VGND VPWR VPWR _191_ sky130_fd_sc_hd__or3_1
XFILLER_12_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_414_ net68 net57 VGND VGND VPWR VPWR _356_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_8_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_800_ clknet_1_0__leaf_clk _002_ _010_ VGND VGND VPWR VPWR tcount\[2\] sky130_fd_sc_hd__dfrtp_2
X_662_ net51 _372_ net20 _076_ VGND VGND VPWR VPWR _222_ sky130_fd_sc_hd__a22o_1
X_731_ net55 net19 _349_ _371_ VGND VGND VPWR VPWR _287_ sky130_fd_sc_hd__a211o_1
XFILLER_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_593_ net71 net59 net51 VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__a21oi_2
XFILLER_6_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput8 net8 VGND VGND VPWR VPWR sine_out[15] sky130_fd_sc_hd__buf_2
X_645_ net41 _063_ _198_ _205_ _369_ VGND VGND VPWR VPWR _206_ sky130_fd_sc_hd__a32o_1
X_576_ _139_ net28 _138_ VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__or3b_1
X_714_ net38 _020_ _096_ _270_ VGND VGND VPWR VPWR _271_ sky130_fd_sc_hd__o31a_1
Xoutput10 net10 VGND VGND VPWR VPWR sine_out[2] sky130_fd_sc_hd__buf_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_430_ net61 net71 VGND VGND VPWR VPWR _372_ sky130_fd_sc_hd__nand2b_4
X_628_ _178_ _179_ _189_ VGND VGND VPWR VPWR _190_ sky130_fd_sc_hd__a21oi_1
X_559_ _344_ _363_ _122_ _121_ _031_ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__o311a_1
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_413_ net70 net56 VGND VGND VPWR VPWR _355_ sky130_fd_sc_hd__and2_1
XFILLER_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_592_ net43 _154_ VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__nand2_1
X_661_ net59 _001_ _036_ net24 VGND VGND VPWR VPWR _221_ sky130_fd_sc_hd__a211o_1
X_730_ _373_ _019_ _075_ _353_ net26 VGND VGND VPWR VPWR _286_ sky130_fd_sc_hd__o221a_1
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_644_ _355_ _361_ net28 VGND VGND VPWR VPWR _205_ sky130_fd_sc_hd__o21a_1
X_575_ net72 net53 net61 net66 VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__and4b_1
XFILLER_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput11 net11 VGND VGND VPWR VPWR sine_out[3] sky130_fd_sc_hd__buf_2
X_713_ _261_ _269_ net26 VGND VGND VPWR VPWR _270_ sky130_fd_sc_hd__a21o_1
Xoutput9 net9 VGND VGND VPWR VPWR sine_out[1] sky130_fd_sc_hd__buf_2
XFILLER_26_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_627_ tcount\[6\] _186_ _188_ _051_ _182_ VGND VGND VPWR VPWR _189_ sky130_fd_sc_hd__a32o_1
X_489_ _000_ _380_ _038_ net47 _032_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__a221oi_1
X_558_ net36 _361_ VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__nand2_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_412_ net57 net63 VGND VGND VPWR VPWR _354_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_591_ net53 net66 _026_ _076_ net22 VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__a32o_1
X_660_ _029_ _042_ _219_ net37 VGND VGND VPWR VPWR _220_ sky130_fd_sc_hd__a22o_1
XFILLER_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_789_ _335_ _336_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__and2_1
Xoutput12 net12 VGND VGND VPWR VPWR sine_out[4] sky130_fd_sc_hd__buf_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_712_ net19 _018_ VGND VGND VPWR VPWR _269_ sky130_fd_sc_hd__nand2_1
XFILLER_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_574_ net52 net66 _363_ VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__or3_1
XFILLER_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_643_ _201_ _203_ _347_ VGND VGND VPWR VPWR _204_ sky130_fd_sc_hd__o21a_1
XFILLER_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_557_ _362_ _390_ _090_ _343_ net44 VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__a221o_1
X_626_ _029_ _049_ _187_ net43 _337_ VGND VGND VPWR VPWR _188_ sky130_fd_sc_hd__a221o_1
X_488_ _347_ _383_ _034_ _053_ VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__a211o_1
XFILLER_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_411_ net55 net62 VGND VGND VPWR VPWR _353_ sky130_fd_sc_hd__and2b_1
X_609_ net29 _170_ _171_ _347_ VGND VGND VPWR VPWR _172_ sky130_fd_sc_hd__o211a_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_24_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_590_ net29 net20 _152_ _348_ VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__a31o_1
X_788_ net34 net43 _128_ tcount\[6\] VGND VGND VPWR VPWR _336_ sky130_fd_sc_hd__a31o_1
XFILLER_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput13 net13 VGND VGND VPWR VPWR sine_out[5] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_11_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_573_ net23 _028_ net20 net52 net42 VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__a221o_1
X_711_ net30 _265_ _268_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__a21bo_1
X_642_ _115_ _202_ net35 VGND VGND VPWR VPWR _203_ sky130_fd_sc_hd__a21oi_1
XFILLER_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_625_ net60 _076_ _364_ VGND VGND VPWR VPWR _187_ sky130_fd_sc_hd__a21bo_1
X_487_ net41 _043_ _044_ _050_ _051_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__o311a_1
X_556_ _385_ _039_ _042_ _348_ VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__a31o_1
XFILLER_8_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_410_ net71 net59 VGND VGND VPWR VPWR _352_ sky130_fd_sc_hd__nand2b_1
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_539_ _026_ _028_ _103_ VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__a21o_1
X_608_ net50 net20 _057_ _372_ net38 VGND VGND VPWR VPWR _171_ sky130_fd_sc_hd__a221o_1
XFILLER_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout70 tcount\[0\] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_2
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_787_ _032_ _334_ VGND VGND VPWR VPWR _335_ sky130_fd_sc_hd__or2_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_572_ _132_ _133_ _135_ _348_ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__a31o_1
X_710_ net30 _258_ _264_ _267_ VGND VGND VPWR VPWR _268_ sky130_fd_sc_hd__or4_1
Xoutput14 net14 VGND VGND VPWR VPWR sine_out[6] sky130_fd_sc_hd__buf_2
X_641_ net24 _351_ _036_ VGND VGND VPWR VPWR _202_ sky130_fd_sc_hd__or3_1
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_486_ _331_ net34 VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__nand2_4
X_624_ net29 _377_ _183_ _185_ net33 VGND VGND VPWR VPWR _186_ sky130_fd_sc_hd__a311o_1
X_555_ net46 _373_ _063_ net35 VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__o211a_1
XFILLER_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_538_ net50 _349_ net26 VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__a21o_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_607_ net24 _367_ _025_ _092_ VGND VGND VPWR VPWR _170_ sky130_fd_sc_hd__o31a_1
X_469_ net59 net65 net71 VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__and3b_1
Xfanout60 net61 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout71 net72 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_4
XFILLER_1_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_786_ net34 _334_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput15 net15 VGND VGND VPWR VPWR sine_out[7] sky130_fd_sc_hd__buf_2
X_571_ net27 _349_ _134_ VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__or3b_1
XFILLER_16_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_640_ net45 _353_ _025_ _361_ net35 VGND VGND VPWR VPWR _201_ sky130_fd_sc_hd__o311a_1
X_769_ net40 net49 _359_ _389_ VGND VGND VPWR VPWR _323_ sky130_fd_sc_hd__a31o_1
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_485_ tcount\[6\] _337_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__nor2_4
X_623_ net28 _380_ _082_ _139_ VGND VGND VPWR VPWR _185_ sky130_fd_sc_hd__nor4_1
XFILLER_12_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_554_ net35 _019_ _041_ _066_ _117_ VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_20_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_468_ net69 net57 net64 VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__or3_1
X_537_ net71 _380_ _101_ net37 VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__a211o_1
X_606_ _051_ _149_ _168_ net30 VGND VGND VPWR VPWR _169_ sky130_fd_sc_hd__a31o_1
X_399_ net71 net65 VGND VGND VPWR VPWR _342_ sky130_fd_sc_hd__nor2_1
XFILLER_4_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout61 tcount\[2\] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_2
Xfanout72 tcount\[0\] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_2
Xfanout50 net54 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_2
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_785_ _129_ _334_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_6_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_570_ net48 _356_ _359_ VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__and3_1
Xoutput16 net16 VGND VGND VPWR VPWR sine_out[8] sky130_fd_sc_hd__buf_2
X_768_ net40 _350_ _134_ VGND VGND VPWR VPWR _322_ sky130_fd_sc_hd__a21oi_1
XFILLER_24_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_22_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_699_ net25 _355_ _106_ VGND VGND VPWR VPWR _257_ sky130_fd_sc_hd__or3_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_622_ net29 _377_ _183_ net33 VGND VGND VPWR VPWR _184_ sky130_fd_sc_hd__a31o_1
X_484_ net27 _048_ _049_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__or3b_1
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_553_ _115_ _116_ net35 VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__a21oi_1
X_398_ net1 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__inv_2
X_467_ _387_ _017_ _030_ _033_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__a2bb2o_1
X_536_ net47 _027_ _072_ VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__and3_1
X_605_ net37 _072_ VGND VGND VPWR VPWR _168_ sky130_fd_sc_hd__or2_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout40 net41 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
Xfanout51 net54 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_4
Xfanout62 net64 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_519_ net51 _021_ _376_ net37 VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_3_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_784_ net43 _128_ VGND VGND VPWR VPWR _334_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_6_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput17 net17 VGND VGND VPWR VPWR sine_out[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_26_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_767_ net27 _320_ VGND VGND VPWR VPWR _321_ sky130_fd_sc_hd__and2_1
XFILLER_30_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_698_ _340_ _066_ _107_ net36 VGND VGND VPWR VPWR _256_ sky130_fd_sc_hd__a31o_1
XFILLER_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_621_ _379_ _064_ VGND VGND VPWR VPWR _183_ sky130_fd_sc_hd__nor2_1
X_483_ net60 _346_ _339_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__a21o_1
X_552_ _351_ _041_ VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__or2_1
XFILLER_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_397_ net31 VGND VGND VPWR VPWR _341_ sky130_fd_sc_hd__inv_2
X_466_ net27 _366_ _020_ _024_ _031_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__o41a_1
X_604_ net39 _042_ _166_ _160_ _032_ VGND VGND VPWR VPWR _167_ sky130_fd_sc_hd__a311o_1
X_535_ _099_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__inv_2
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout41 net44 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
Xfanout52 net54 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_2
Xfanout63 net64 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_4
Xfanout30 net32 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_449_ net24 _390_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__nand2_1
X_518_ net37 _082_ VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__nor2_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_783_ _090_ _128_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__nor2_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_766_ net49 _359_ _076_ net58 VGND VGND VPWR VPWR _320_ sky130_fd_sc_hd__a22o_1
X_697_ net45 _197_ _254_ VGND VGND VPWR VPWR _255_ sky130_fd_sc_hd__a21o_1
XFILLER_7_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_620_ net28 _060_ _161_ _180_ _181_ VGND VGND VPWR VPWR _182_ sky130_fd_sc_hd__o32ai_1
XFILLER_21_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_551_ net45 net19 _353_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_749_ _016_ _023_ _063_ net42 VGND VGND VPWR VPWR _304_ sky130_fd_sc_hd__a31o_1
X_482_ _359_ net18 VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_3_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_465_ tcount\[6\] net33 VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__nand2_4
X_396_ net64 VGND VGND VPWR VPWR _340_ sky130_fd_sc_hd__inv_2
X_603_ _344_ _082_ VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__or2_1
X_534_ _032_ _088_ _094_ _098_ net30 VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__o311a_1
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout31 net32 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
Xfanout53 net54 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout42 net43 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
Xfanout64 tcount\[1\] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout20 _037_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_4
X_448_ net72 net66 net60 VGND VGND VPWR VPWR _390_ sky130_fd_sc_hd__a21bo_2
X_517_ net53 net60 net72 VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_0_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_782_ net32 _332_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__and2_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_765_ net34 _316_ _317_ _318_ VGND VGND VPWR VPWR _319_ sky130_fd_sc_hd__a31o_1
X_696_ net25 _390_ net36 VGND VGND VPWR VPWR _254_ sky130_fd_sc_hd__a21o_1
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_550_ net46 _111_ _105_ VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__a21o_1
X_481_ net45 _351_ _045_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__nor3_1
X_748_ _161_ _294_ _179_ VGND VGND VPWR VPWR _303_ sky130_fd_sc_hd__or3b_1
X_679_ net52 _027_ _072_ _237_ VGND VGND VPWR VPWR _238_ sky130_fd_sc_hd__a31o_1
X_464_ _331_ _337_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__nor2_4
X_533_ net29 _095_ _097_ _052_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__a211o_1
X_602_ _151_ _153_ _163_ _032_ net30 VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__o221a_1
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_395_ net51 VGND VGND VPWR VPWR _339_ sky130_fd_sc_hd__inv_2
Xfanout32 tcount\[7\] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_2
Xfanout43 net44 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
Xfanout54 tcount\[3\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
Xfanout21 _389_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_4
Xfanout65 net66 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_447_ tcount\[6\] net33 VGND VGND VPWR VPWR _389_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_516_ net65 _351_ _364_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__a21o_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_781_ net31 _330_ _333_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__a21oi_1
XFILLER_27_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_7_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_764_ _337_ net40 _091_ _331_ VGND VGND VPWR VPWR _318_ sky130_fd_sc_hd__a31o_1
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_695_ net27 net18 _241_ VGND VGND VPWR VPWR _253_ sky130_fd_sc_hd__or3_1
XFILLER_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_480_ net48 _045_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_14_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_678_ net29 _379_ _380_ VGND VGND VPWR VPWR _237_ sky130_fd_sc_hd__or3_1
X_747_ _301_ _302_ net30 _298_ VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__o2bb2a_1
XFILLER_7_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_601_ _052_ _150_ _159_ VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__o21a_1
XFILLER_5_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_463_ _027_ _029_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__nand2_1
X_532_ _344_ _026_ _039_ net37 VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__o211a_1
X_394_ net38 VGND VGND VPWR VPWR _338_ sky130_fd_sc_hd__inv_2
Xfanout33 net34 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_4
Xfanout44 tcount\[4\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout22 _360_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
Xfanout55 net56 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
X_446_ tcount\[6\] net33 VGND VGND VPWR VPWR _388_ sky130_fd_sc_hd__nor2_4
Xfanout66 tcount\[1\] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_2
XFILLER_13_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_515_ net36 _062_ _078_ _079_ VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_23_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_429_ net55 net70 VGND VGND VPWR VPWR _371_ sky130_fd_sc_hd__and2b_2
X_780_ _330_ _332_ net31 VGND VGND VPWR VPWR _333_ sky130_fd_sc_hd__a21oi_1
Xinput1 rst VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_763_ _349_ _363_ _134_ net40 VGND VGND VPWR VPWR _317_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_17_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_694_ net36 _047_ _251_ _250_ VGND VGND VPWR VPWR _252_ sky130_fd_sc_hd__o31ai_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_677_ _031_ _233_ _235_ _232_ _347_ VGND VGND VPWR VPWR _236_ sky130_fd_sc_hd__a32o_1
X_746_ net30 _289_ _292_ VGND VGND VPWR VPWR _302_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_393_ net34 VGND VGND VPWR VPWR _337_ sky130_fd_sc_hd__inv_2
XFILLER_27_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_462_ net25 _354_ net41 VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__a21oi_2
X_600_ net37 _162_ _160_ VGND VGND VPWR VPWR _163_ sky130_fd_sc_hd__a21oi_1
X_531_ _357_ _371_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__nor2_1
X_729_ net26 _283_ _284_ _347_ VGND VGND VPWR VPWR _285_ sky130_fd_sc_hd__o211ai_1
Xfanout34 tcount\[5\] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_4
Xfanout23 _346_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout67 net70 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_4
Xfanout45 net46 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_514_ _051_ _068_ _073_ _031_ net26 VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__a221o_1
Xfanout56 tcount\[2\] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
X_445_ net22 _361_ _385_ _386_ VGND VGND VPWR VPWR _387_ sky130_fd_sc_hd__o22a_1
X_428_ net42 _369_ VGND VGND VPWR VPWR _370_ sky130_fd_sc_hd__nand2_1
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_762_ net68 _384_ _134_ net40 VGND VGND VPWR VPWR _316_ sky130_fd_sc_hd__a211o_1
XFILLER_24_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_693_ net45 _345_ _026_ VGND VGND VPWR VPWR _251_ sky130_fd_sc_hd__and3_1
XFILLER_30_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_676_ _345_ _107_ _234_ net27 VGND VGND VPWR VPWR _235_ sky130_fd_sc_hd__a211o_1
X_745_ _295_ _299_ _300_ net21 VGND VGND VPWR VPWR _301_ sky130_fd_sc_hd__a31o_1
X_392_ tcount\[6\] VGND VGND VPWR VPWR _331_ sky130_fd_sc_hd__inv_2
XFILLER_27_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_530_ net50 _340_ _363_ _380_ _344_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__a311o_1
X_461_ net50 _353_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__nor2_1
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_728_ _343_ _374_ net41 VGND VGND VPWR VPWR _284_ sky130_fd_sc_hd__a21o_1
X_659_ net50 _352_ _022_ _358_ _340_ VGND VGND VPWR VPWR _219_ sky130_fd_sc_hd__a32o_1
Xfanout57 tcount\[2\] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_4
Xfanout68 net70 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout46 net49 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout35 net39 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
Xfanout24 net25 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
X_444_ net69 net44 VGND VGND VPWR VPWR _386_ sky130_fd_sc_hd__nor2_1
X_513_ _075_ _077_ _348_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__a21oi_1
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_427_ net60 net23 _368_ net24 VGND VGND VPWR VPWR _369_ sky130_fd_sc_hd__o211ai_2
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_761_ net31 _306_ _313_ _315_ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__a31o_1
XFILLER_21_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_692_ net27 net62 _363_ _018_ _249_ VGND VGND VPWR VPWR _250_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_22_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_675_ net58 _039_ VGND VGND VPWR VPWR _234_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_744_ net35 net25 _026_ VGND VGND VPWR VPWR _300_ sky130_fd_sc_hd__or3_1
XFILLER_27_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_460_ net64 _026_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__or2_1
X_391_ net72 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_727_ net50 _342_ _351_ _367_ _357_ VGND VGND VPWR VPWR _283_ sky130_fd_sc_hd__o41a_1
X_658_ _032_ _215_ _217_ VGND VGND VPWR VPWR _218_ sky130_fd_sc_hd__or3_1
X_589_ _345_ _028_ VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__nand2_1
Xfanout47 net49 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
Xfanout58 tcount\[2\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout69 net70 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_1
Xfanout36 net39 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout25 _339_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_4
X_443_ net40 _384_ VGND VGND VPWR VPWR _385_ sky130_fd_sc_hd__nor2_1
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_512_ net22 _076_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__nand2_1
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_426_ net72 net66 net60 VGND VGND VPWR VPWR _368_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_1_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_27_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_409_ net67 net55 VGND VGND VPWR VPWR _351_ sky130_fd_sc_hd__and2b_2
XFILLER_24_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_760_ _306_ _314_ net31 VGND VGND VPWR VPWR _315_ sky130_fd_sc_hd__a21oi_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_691_ net26 net45 _070_ VGND VGND VPWR VPWR _249_ sky130_fd_sc_hd__or3_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_674_ net25 _072_ _074_ _354_ net41 VGND VGND VPWR VPWR _233_ sky130_fd_sc_hd__a221o_1
X_743_ net35 _069_ _092_ VGND VGND VPWR VPWR _299_ sky130_fd_sc_hd__or3_1
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_14_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_726_ net32 _281_ _282_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__a21o_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_657_ net26 _202_ _216_ VGND VGND VPWR VPWR _217_ sky130_fd_sc_hd__and3_1
XFILLER_4_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_588_ _364_ _373_ _092_ net38 VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__o211a_1
Xfanout48 net49 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_2
Xfanout59 net61 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_2
Xfanout37 net38 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
Xfanout26 net29 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_2
X_442_ net48 net57 net63 VGND VGND VPWR VPWR _384_ sky130_fd_sc_hd__and3b_1
XFILLER_1_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_511_ net71 net65 net51 VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__o21ba_4
X_709_ _250_ _266_ net21 VGND VGND VPWR VPWR _267_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_425_ net65 net59 VGND VGND VPWR VPWR _367_ sky130_fd_sc_hd__and2b_2
XFILLER_27_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_408_ net58 net64 VGND VGND VPWR VPWR _350_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_2_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_690_ net31 _247_ _248_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__o21ai_1
XFILLER_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_673_ _366_ _231_ _230_ _385_ VGND VGND VPWR VPWR _232_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_742_ _289_ _292_ _297_ VGND VGND VPWR VPWR _298_ sky130_fd_sc_hd__and3_1
X_587_ net37 _363_ _367_ _149_ VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__o31a_1
X_725_ net21 _271_ _278_ _341_ VGND VGND VPWR VPWR _282_ sky130_fd_sc_hd__o211a_1
X_656_ net20 _076_ VGND VGND VPWR VPWR _216_ sky130_fd_sc_hd__nand2_1
Xfanout49 net54 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_2
Xfanout27 net28 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
Xfanout38 net39 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
X_441_ _365_ _370_ _382_ VGND VGND VPWR VPWR _383_ sky130_fd_sc_hd__o21ai_1
X_510_ net56 net19 _364_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__a21o_1
X_639_ net41 _048_ _058_ _199_ _031_ VGND VGND VPWR VPWR _200_ sky130_fd_sc_hd__o311a_1
X_708_ net67 _018_ _251_ net36 VGND VGND VPWR VPWR _266_ sky130_fd_sc_hd__a211o_1
XFILLER_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_424_ net59 net23 VGND VGND VPWR VPWR _366_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_407_ net55 net62 VGND VGND VPWR VPWR _349_ sky130_fd_sc_hd__nor2_2
XFILLER_15_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_672_ net36 _066_ VGND VGND VPWR VPWR _231_ sky130_fd_sc_hd__nand2_1
X_741_ _295_ _296_ net21 VGND VGND VPWR VPWR _297_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_724_ _278_ _280_ VGND VGND VPWR VPWR _281_ sky130_fd_sc_hd__nand2_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_586_ net59 _076_ _126_ _067_ VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__a211o_1
X_655_ net50 _366_ _377_ net38 VGND VGND VPWR VPWR _215_ sky130_fd_sc_hd__o211a_1
X_440_ net42 _378_ _379_ _380_ VGND VGND VPWR VPWR _382_ sky130_fd_sc_hd__or4_1
Xfanout28 net29 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_2
Xfanout39 net44 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlymetal6s2s_1
X_638_ _354_ _356_ _198_ _067_ net28 VGND VGND VPWR VPWR _199_ sky130_fd_sc_hd__a311o_1
X_569_ net47 _045_ _106_ VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__or3_1
X_707_ _388_ _252_ _258_ _264_ VGND VGND VPWR VPWR _265_ sky130_fd_sc_hd__a211o_1
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_423_ _000_ _339_ _360_ VGND VGND VPWR VPWR _365_ sky130_fd_sc_hd__nor3_1
XFILLER_10_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_406_ tcount\[6\] _337_ VGND VGND VPWR VPWR _348_ sky130_fd_sc_hd__nand2_2
XFILLER_18_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_671_ _344_ _364_ VGND VGND VPWR VPWR _230_ sky130_fd_sc_hd__or2_1
XFILLER_11_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_740_ net36 _351_ _384_ _260_ VGND VGND VPWR VPWR _296_ sky130_fd_sc_hd__or4_1
XFILLER_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_654_ _212_ _213_ _388_ VGND VGND VPWR VPWR _214_ sky130_fd_sc_hd__o21ai_1
X_585_ _124_ _125_ _148_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__o21ba_1
X_723_ _270_ _279_ net21 VGND VGND VPWR VPWR _280_ sky130_fd_sc_hd__a21o_1
XFILLER_1_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout29 _338_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_2
X_637_ net68 _354_ _359_ _069_ net48 VGND VGND VPWR VPWR _198_ sky130_fd_sc_hd__a221o_1
X_706_ _031_ _253_ _255_ _263_ VGND VGND VPWR VPWR _264_ sky130_fd_sc_hd__a31o_1
X_499_ net52 net60 VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__nor2_1
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_568_ _022_ _028_ _040_ _057_ net42 VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__a221o_1
X_422_ net70 net56 net49 VGND VGND VPWR VPWR _364_ sky130_fd_sc_hd__o21ai_4
XFILLER_6_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_405_ _331_ net34 VGND VGND VPWR VPWR _347_ sky130_fd_sc_hd__nor2_4
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_20_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_670_ _214_ _225_ _229_ _341_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__a22oi_1
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_799_ clknet_1_0__leaf_clk net19 _009_ VGND VGND VPWR VPWR tcount\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_584_ _130_ _141_ _147_ _136_ VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__and4bb_1
X_653_ _087_ _112_ net26 VGND VGND VPWR VPWR _213_ sky130_fd_sc_hd__o21a_1
X_722_ _018_ _057_ _096_ net38 VGND VGND VPWR VPWR _279_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_9_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout19 _001_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XFILLER_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_498_ net53 _360_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__nand2_2
X_705_ net27 _074_ _259_ _262_ _347_ VGND VGND VPWR VPWR _263_ sky130_fd_sc_hd__o311a_1
X_636_ net68 net22 _022_ _356_ VGND VGND VPWR VPWR _197_ sky130_fd_sc_hd__o211a_1
X_567_ _040_ _057_ net37 VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_421_ net68 net57 VGND VGND VPWR VPWR _363_ sky130_fd_sc_hd__nor2_2
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_619_ net72 net52 net60 net43 VGND VGND VPWR VPWR _181_ sky130_fd_sc_hd__a31o_1
XFILLER_14_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_404_ net23 VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_22_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_798_ clknet_1_0__leaf_clk _000_ _008_ VGND VGND VPWR VPWR tcount\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_583_ _143_ _144_ _146_ _052_ VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__a31o_1
X_721_ _131_ _272_ _274_ _277_ VGND VGND VPWR VPWR _278_ sky130_fd_sc_hd__o211a_1
X_652_ net66 _156_ _103_ VGND VGND VPWR VPWR _212_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_635_ _193_ _195_ net21 VGND VGND VPWR VPWR _196_ sky130_fd_sc_hd__a21oi_1
X_566_ _370_ _126_ _127_ _129_ _388_ VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__o221a_1
X_704_ net48 _354_ _356_ _260_ net41 VGND VGND VPWR VPWR _262_ sky130_fd_sc_hd__a311o_1
X_497_ _347_ _055_ _061_ _051_ _054_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__a221o_1
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_420_ _361_ VGND VGND VPWR VPWR _362_ sky130_fd_sc_hd__inv_2
X_618_ net60 net23 _156_ VGND VGND VPWR VPWR _180_ sky130_fd_sc_hd__o21a_1
X_549_ _096_ _112_ net35 VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__o21ai_1
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_403_ net71 net65 VGND VGND VPWR VPWR _346_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_19_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_797_ net1 VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__inv_2
XFILLER_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_651_ _208_ _211_ _341_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__mux2_1
X_582_ net28 net19 _364_ VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__or3_1
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_720_ net26 _025_ _275_ _276_ _032_ VGND VGND VPWR VPWR _277_ sky130_fd_sc_hd__a311o_1
XFILLER_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_565_ net43 _128_ VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__or2_1
X_634_ net18 _194_ VGND VGND VPWR VPWR _195_ sky130_fd_sc_hd__or2_1
X_496_ _372_ _040_ _057_ _060_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__a31oi_1
X_703_ _342_ _026_ net50 VGND VGND VPWR VPWR _261_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_617_ _345_ _064_ VGND VGND VPWR VPWR _179_ sky130_fd_sc_hd__nand2_1
X_479_ net57 net63 net68 VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__nor3b_4
X_548_ net20 _111_ net46 VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__a21oi_1
XFILLER_25_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_402_ net68 net63 VGND VGND VPWR VPWR _345_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_19_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap18 _047_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_16_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_796_ net1 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__inv_2
X_650_ _200_ _204_ _207_ _210_ VGND VGND VPWR VPWR _211_ sky130_fd_sc_hd__and4bb_1
X_779_ tcount\[6\] net33 _325_ VGND VGND VPWR VPWR _332_ sky130_fd_sc_hd__or3_1
X_581_ net43 net47 VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_564_ net72 net52 net60 tcount\[1\] VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__and4_1
X_633_ net47 _343_ _037_ net40 VGND VGND VPWR VPWR _194_ sky130_fd_sc_hd__a31o_1
X_495_ _339_ net22 _022_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__and3_1
XFILLER_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_702_ net55 net46 net67 VGND VGND VPWR VPWR _260_ sky130_fd_sc_hd__and3b_1
XFILLER_5_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_616_ net28 _176_ _177_ _388_ VGND VGND VPWR VPWR _178_ sky130_fd_sc_hd__o211a_1
X_478_ net48 net63 _363_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__and3_1
X_547_ net22 _372_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__nand2_1
XFILLER_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_401_ net72 net65 VGND VGND VPWR VPWR _344_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_19_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_795_ net1 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__inv_2
X_580_ _343_ _350_ _359_ net47 net27 VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_4_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_778_ _388_ _145_ _325_ _284_ _031_ VGND VGND VPWR VPWR _330_ sky130_fd_sc_hd__a32oi_2
XPHY_EDGE_ROW_13_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_632_ _044_ _192_ net40 VGND VGND VPWR VPWR _193_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_563_ net52 _072_ VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__nor2_1
X_701_ _346_ _065_ _371_ VGND VGND VPWR VPWR _259_ sky130_fd_sc_hd__a21oi_1
X_494_ net25 net22 VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__and2_1
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_615_ net25 net22 _386_ VGND VGND VPWR VPWR _177_ sky130_fd_sc_hd__or3b_1
X_477_ net19 _040_ _038_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__a21oi_1
XFILLER_14_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_546_ net30 _080_ _085_ _100_ _110_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__o32a_1
X_400_ net69 net64 VGND VGND VPWR VPWR _343_ sky130_fd_sc_hd__or2_1
XFILLER_17_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_529_ _069_ _092_ _093_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__o21a_1
XFILLER_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_794_ net1 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__inv_2
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_777_ _329_ _341_ _328_ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__mux2_1
X_700_ _249_ _256_ _257_ _052_ VGND VGND VPWR VPWR _258_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_631_ net69 net22 _361_ _089_ VGND VGND VPWR VPWR _192_ sky130_fd_sc_hd__o22a_1
X_493_ _349_ _042_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__nor2_1
X_562_ _357_ _358_ _045_ VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_614_ _027_ _107_ VGND VGND VPWR VPWR _176_ sky130_fd_sc_hd__nor2_1
X_476_ net51 _372_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__nand2_2
X_545_ _388_ _102_ _104_ _109_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_1_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_459_ net67 net55 VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__xor2_4
X_528_ net24 _351_ _021_ net38 VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__o31a_1
XFILLER_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_793_ net1 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__inv_2
XFILLER_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_776_ net33 _325_ net31 VGND VGND VPWR VPWR _329_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_630_ _341_ _190_ _191_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__o21ai_1
XFILLER_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_561_ _388_ _113_ _114_ _123_ VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__a31o_1
X_492_ net56 net19 VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__nand2_1
XFILLER_5_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_759_ _184_ _311_ _309_ VGND VGND VPWR VPWR _314_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_613_ _164_ _165_ _174_ _175_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__o2bb2a_1
X_544_ _101_ _105_ _108_ _347_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__o211a_1
X_475_ net67 net62 net45 VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_28_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_527_ _045_ _091_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__or2_1
XFILLER_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_458_ _351_ _371_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_30_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_792_ net1 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__inv_2
XFILLER_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_775_ _347_ _327_ VGND VGND VPWR VPWR _328_ sky130_fd_sc_hd__or2_1
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_491_ _342_ _390_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__nor2_1
X_560_ _052_ _118_ _119_ _120_ net30 VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__o221ai_1
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_689_ _240_ _244_ _341_ _236_ VGND VGND VPWR VPWR _248_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_758_ _309_ _312_ VGND VGND VPWR VPWR _313_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_17_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_543_ _375_ _022_ _065_ _106_ VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__a31o_1
X_474_ _375_ _039_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__nand2_1
X_612_ _169_ _172_ _167_ VGND VGND VPWR VPWR _175_ sky130_fd_sc_hd__or3b_1
XFILLER_26_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_526_ net68 net57 net63 net48 VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__a31o_1
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_457_ _375_ _022_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__nor2_1
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_509_ net57 net19 _364_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_791_ net1 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_774_ _051_ _183_ _284_ _145_ VGND VGND VPWR VPWR _327_ sky130_fd_sc_hd__a22o_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_490_ _345_ _018_ _025_ _036_ net50 VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__a32o_1
X_757_ net29 _377_ _310_ _311_ net33 VGND VGND VPWR VPWR _312_ sky130_fd_sc_hd__a311o_1
X_688_ _240_ _246_ _236_ VGND VGND VPWR VPWR _247_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_542_ _375_ _065_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__nand2_1
X_611_ net42 _173_ _155_ _388_ VGND VGND VPWR VPWR _174_ sky130_fd_sc_hd__o211a_1
X_473_ net46 net64 VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__nand2_1
XFILLER_26_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_525_ net47 _089_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__nor2_1
X_456_ net52 _355_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_439_ net24 _367_ VGND VGND VPWR VPWR _381_ sky130_fd_sc_hd__nand2_1
X_508_ net25 _072_ _071_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_30_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_790_ net32 _335_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_12_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_773_ _341_ _326_ _324_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__mux2_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_687_ _242_ _245_ net34 VGND VGND VPWR VPWR _246_ sky130_fd_sc_hd__a21o_1
XFILLER_18_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_756_ net24 _367_ _036_ _086_ net39 VGND VGND VPWR VPWR _311_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_5_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_472_ _390_ _035_ _037_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__and3_1
X_610_ _000_ _376_ _065_ VGND VGND VPWR VPWR _173_ sky130_fd_sc_hd__o21a_1
X_541_ _000_ net66 net28 VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__a21o_1
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_739_ net20 _111_ _293_ _294_ VGND VGND VPWR VPWR _295_ sky130_fd_sc_hd__a31o_1
X_524_ net69 net58 net63 VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__and3_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_455_ net62 net67 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_2_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_438_ net51 net65 net61 VGND VGND VPWR VPWR _380_ sky130_fd_sc_hd__nor3b_2
X_507_ net62 _026_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__nand2_2
XFILLER_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_772_ net31 _325_ VGND VGND VPWR VPWR _326_ sky130_fd_sc_hd__and2_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_755_ _368_ net20 net53 VGND VGND VPWR VPWR _310_ sky130_fd_sc_hd__a21o_1
X_686_ _385_ _142_ VGND VGND VPWR VPWR _245_ sky130_fd_sc_hd__nand2_1
XFILLER_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_471_ _390_ net20 VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__nand2_1
X_540_ _385_ _066_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__nand2_1
X_738_ net27 _384_ VGND VGND VPWR VPWR _294_ sky130_fd_sc_hd__or2_1
X_669_ _052_ _220_ _226_ _227_ _228_ VGND VGND VPWR VPWR _229_ sky130_fd_sc_hd__o2111a_1
XFILLER_26_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_523_ _349_ _355_ _364_ _086_ net29 VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__o311a_1
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_454_ net66 net71 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_18_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_437_ net72 net52 net66 VGND VGND VPWR VPWR _379_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_15_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_506_ net45 _070_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_771_ net43 _179_ VGND VGND VPWR VPWR _325_ sky130_fd_sc_hd__or2_1
XFILLER_3_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_685_ _242_ _243_ net34 VGND VGND VPWR VPWR _244_ sky130_fd_sc_hd__a21o_1
X_754_ net33 _307_ _308_ tcount\[6\] VGND VGND VPWR VPWR _309_ sky130_fd_sc_hd__a31oi_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_599_ net61 _076_ _161_ _067_ VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__a211o_1
X_668_ net26 _381_ _142_ _212_ net21 VGND VGND VPWR VPWR _228_ sky130_fd_sc_hd__a311o_1
X_470_ net59 net65 net71 VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__nand3b_2
X_737_ _372_ _076_ VGND VGND VPWR VPWR _293_ sky130_fd_sc_hd__nand2_1
XFILLER_17_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_522_ _349_ _364_ VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__nor2_1
X_453_ net19 _019_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__nor2_1
Xoutput2 net2 VGND VGND VPWR VPWR sine_out[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_18_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_436_ _371_ _377_ VGND VGND VPWR VPWR _378_ sky130_fd_sc_hd__nor2_1
X_505_ net55 net62 net67 VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__o21bai_1
XFILLER_22_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_25_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_419_ net68 net63 net47 VGND VGND VPWR VPWR _361_ sky130_fd_sc_hd__o21ai_4
X_770_ _052_ _321_ _322_ _323_ _319_ VGND VGND VPWR VPWR _324_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_684_ net40 _349_ _363_ _384_ VGND VGND VPWR VPWR _243_ sky130_fd_sc_hd__or4_1
X_753_ net42 _065_ VGND VGND VPWR VPWR _308_ sky130_fd_sc_hd__nand2_1
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_12_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_805_ clknet_1_1__leaf_clk _007_ _015_ VGND VGND VPWR VPWR tcount\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_736_ net38 _290_ _291_ _052_ VGND VGND VPWR VPWR _292_ sky130_fd_sc_hd__a211o_1
XFILLER_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_598_ _368_ net20 net25 VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__a21oi_1
X_667_ _347_ _223_ VGND VGND VPWR VPWR _227_ sky130_fd_sc_hd__nand2_1
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_452_ net56 net62 net46 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__o21bai_2
X_521_ net51 _360_ _021_ VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__or3_1
Xoutput3 net3 VGND VGND VPWR VPWR sine_out[10] sky130_fd_sc_hd__buf_2
X_719_ _361_ _367_ _019_ net23 net35 VGND VGND VPWR VPWR _276_ sky130_fd_sc_hd__o221a_1
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_435_ net59 net23 _353_ net24 VGND VGND VPWR VPWR _377_ sky130_fd_sc_hd__a211o_1
X_504_ net56 net62 net67 VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__o21ba_1
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_0_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_418_ net57 net63 VGND VGND VPWR VPWR _360_ sky130_fd_sc_hd__xnor2_4
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_683_ _059_ _241_ net40 VGND VGND VPWR VPWR _242_ sky130_fd_sc_hd__o21ai_1
X_752_ _360_ _372_ _082_ net42 VGND VGND VPWR VPWR _307_ sky130_fd_sc_hd__a211o_1
XFILLER_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_804_ clknet_1_1__leaf_clk _006_ _014_ VGND VGND VPWR VPWR tcount\[6\] sky130_fd_sc_hd__dfrtp_4
X_735_ _001_ _023_ _129_ VGND VGND VPWR VPWR _291_ sky130_fd_sc_hd__a21oi_1
X_597_ net24 _045_ _056_ _083_ VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__o31a_1
X_666_ _215_ _217_ _031_ VGND VGND VPWR VPWR _226_ sky130_fd_sc_hd__o21ai_1
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_520_ _081_ _083_ _084_ net21 VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__a211oi_1
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput4 net4 VGND VGND VPWR VPWR sine_out[11] sky130_fd_sc_hd__buf_2
X_649_ _193_ _209_ _389_ VGND VGND VPWR VPWR _210_ sky130_fd_sc_hd__a21o_1
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_451_ net55 net62 net45 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__o21ba_2
X_718_ net46 net23 VGND VGND VPWR VPWR _275_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_24_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_434_ net48 _354_ VGND VGND VPWR VPWR _376_ sky130_fd_sc_hd__nand2_1
X_503_ net67 net46 net22 _067_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_21_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_417_ net57 net63 VGND VGND VPWR VPWR _359_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_751_ net33 _303_ _304_ _305_ _331_ VGND VGND VPWR VPWR _306_ sky130_fd_sc_hd__a311o_1
XFILLER_18_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_682_ _045_ _069_ net48 VGND VGND VPWR VPWR _241_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_803_ clknet_1_1__leaf_clk _005_ _013_ VGND VGND VPWR VPWR tcount\[5\] sky130_fd_sc_hd__dfrtp_1
X_596_ _155_ _158_ net21 VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__a21o_1
X_665_ net30 _218_ _224_ VGND VGND VPWR VPWR _225_ sky130_fd_sc_hd__and3_1
X_734_ _372_ _028_ VGND VGND VPWR VPWR _290_ sky130_fd_sc_hd__nand2_1
Xoutput5 net5 VGND VGND VPWR VPWR sine_out[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_27_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_450_ net42 _375_ _016_ net21 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__a31o_1
X_648_ net68 _018_ _194_ VGND VGND VPWR VPWR _209_ sky130_fd_sc_hd__a21o_1
X_579_ _026_ _040_ _076_ net41 VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__a211o_1
XFILLER_16_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_717_ net37 _138_ _142_ _273_ _052_ VGND VGND VPWR VPWR _274_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_24_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_433_ net47 net58 VGND VGND VPWR VPWR _375_ sky130_fd_sc_hd__nand2_1
X_502_ _345_ _065_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__nor2_2
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_416_ net61 net51 VGND VGND VPWR VPWR _358_ sky130_fd_sc_hd__nand2b_1
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_750_ _374_ _090_ _035_ _337_ net43 VGND VGND VPWR VPWR _305_ sky130_fd_sc_hd__o2111a_1
X_681_ _331_ _238_ _239_ _388_ VGND VGND VPWR VPWR _240_ sky130_fd_sc_hd__a31o_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_802_ clknet_1_1__leaf_clk _004_ _012_ VGND VGND VPWR VPWR tcount\[4\] sky130_fd_sc_hd__dfrtp_1
X_595_ _023_ _063_ _157_ net42 VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__a31o_1
XFILLER_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_733_ _032_ _286_ _288_ _285_ VGND VGND VPWR VPWR _289_ sky130_fd_sc_hd__o31a_1
X_664_ _051_ _220_ _223_ _348_ VGND VGND VPWR VPWR _224_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput6 net6 VGND VGND VPWR VPWR sine_out[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_27_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_647_ _196_ _200_ _204_ _207_ VGND VGND VPWR VPWR _208_ sky130_fd_sc_hd__or4b_1
X_716_ _355_ _364_ _069_ net50 net28 VGND VGND VPWR VPWR _273_ sky130_fd_sc_hd__o221a_1
X_578_ net55 _041_ VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__or2_2
.ends

